`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/01/2025 10:20:40 PM
// Design Name: 
// Module Name: AXI4L_SLV_IF_64AR
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AXI4L_SLV_IF_64AR # (
		// Width of S_AXI data bus
		parameter integer C_S_AXI_DATA_WIDTH	= 32,
		// Width of S_AXI address bus
		parameter integer C_S_AXI_ADDR_WIDTH	= 10
	)
	(
    // ==================================================================== //
    //  AXI4-Lite Slave Interface Pins                                      //
    // ==================================================================== //
        // General
		input wire                              S_AXI_ACLK,     // AXI CLK
		input wire                              S_AXI_ARESETN,  // AXI RESET (Active Low)

        // Write Address Channel
		input wire [C_S_AXI_ADDR_WIDTH-1:0]     S_AXI_AWADDR,   // Write Address (Issued by Master, Accepted by Slave)
		input wire [2:0]                        S_AXI_AWPROT,   // Write Channel Protection Type
		input wire                              S_AXI_AWVALID,  // Write Address Valid
		output wire                             S_AXI_AWREADY,  // Write Address Ready

        // Write Data Channel
		input wire [C_S_AXI_DATA_WIDTH-1:0]     S_AXI_WDATA,    // Write Data (Issued by Master, Accepted By Slave)   
		input wire [(C_S_AXI_DATA_WIDTH/8)-1:0] S_AXI_WSTRB,    // Write Strobe (Indicates which Byte lanes hold valid data. One Write Strobe bit for Each Eight bits of the Write Data bus)
		input wire                              S_AXI_WVALID,   // Write Valid
		output wire                             S_AXI_WREADY,   // Write Ready

        // Write Response Channel
		output wire [1:0]                       S_AXI_BRESP,    // Write Response
		output wire                             S_AXI_BVALID,   // Write Response Valid           
		input wire                              S_AXI_BREADY,   // Write Response Ready
		
        // Read Address Channel
		input wire [C_S_AXI_ADDR_WIDTH-1:0]     S_AXI_ARADDR,   // Read Address (Issued by Master, Accepted by Slave)
		input wire [2:0]                        S_AXI_ARPROT,   // Read Channel Protection Type
		input wire                              S_AXI_ARVALID,  // Read Address Valid
		output wire                             S_AXI_ARREADY,  // Read Address Ready

        // Read Data Channel
		output wire [C_S_AXI_DATA_WIDTH-1:0]    S_AXI_RDATA,    // Read Data (Issued by Slave, Accepted by Master)
		output wire [1:0]                       S_AXI_RRESP,    // Read Response
		output wire                             S_AXI_RVALID,   // Read Valid
		input wire                              S_AXI_RREADY,   // Read Ready

    // ==================================================================== //
    //  User Custom I/O Pins                                                //
    // ==================================================================== //
        // Add User Input Pins  (# User Guide : Uncomment Pins to Use)
        // input wire [31:0]                       i_reg_64bit_1th_hi,          // Match to 'slv_reg0'
        // input wire [31:0]                       i_reg_64bit_1th_lo,          // Match to 'slv_reg1'
        // input wire [31:0]                       i_reg_64bit_2th_hi,
        // input wire [31:0]                       i_reg_64bit_2th_lo,
        // input wire [31:0]                       i_reg_64bit_3th_hi,
        // input wire [31:0]                       i_reg_64bit_3th_lo,
        // input wire [31:0]                       i_reg_64bit_4th_hi,
        // input wire [31:0]                       i_reg_64bit_4th_lo,
        // input wire [31:0]                       i_reg_64bit_5th_hi,
        // input wire [31:0]                       i_reg_64bit_5th_lo,
        // input wire [31:0]                       i_reg_64bit_6th_hi,
        // input wire [31:0]                       i_reg_64bit_6th_lo,
        // input wire [31:0]                       i_reg_64bit_7th_hi,
        // input wire [31:0]                       i_reg_64bit_7th_lo,
        // input wire [31:0]                       i_reg_64bit_8th_hi,
        // input wire [31:0]                       i_reg_64bit_8th_lo,
        // input wire [31:0]                       i_reg_64bit_9th_hi,
        // input wire [31:0]                       i_reg_64bit_9th_lo,
        // input wire [31:0]                       i_reg_64bit_10th_hi,
        // input wire [31:0]                       i_reg_64bit_10th_lo,
        // input wire [31:0]                       i_reg_64bit_11th_hi,
        // input wire [31:0]                       i_reg_64bit_11th_lo,
        // input wire [31:0]                       i_reg_64bit_12th_hi,
        // input wire [31:0]                       i_reg_64bit_12th_lo,
        // input wire [31:0]                       i_reg_64bit_13th_hi,
        // input wire [31:0]                       i_reg_64bit_13th_lo,
        // input wire [31:0]                       i_reg_64bit_14th_hi,
        // input wire [31:0]                       i_reg_64bit_14th_lo,
        // input wire [31:0]                       i_reg_64bit_15th_hi,
        // input wire [31:0]                       i_reg_64bit_15th_lo,
        // input wire [31:0]                       i_reg_64bit_16th_hi,
        // input wire [31:0]                       i_reg_64bit_16th_lo,
        // input wire [31:0]                       i_reg_64bit_17th_hi,
        // input wire [31:0]                       i_reg_64bit_17th_lo,
        // input wire [31:0]                       i_reg_64bit_18th_hi,
        // input wire [31:0]                       i_reg_64bit_18th_lo,
        // input wire [31:0]                       i_reg_64bit_19th_hi,
        // input wire [31:0]                       i_reg_64bit_19th_lo,
        // input wire [31:0]                       i_reg_64bit_20th_hi,
        // input wire [31:0]                       i_reg_64bit_20th_lo,
        // input wire [31:0]                       i_reg_64bit_21th_hi,
        // input wire [31:0]                       i_reg_64bit_21th_lo,
        // input wire [31:0]                       i_reg_64bit_22th_hi,
        // input wire [31:0]                       i_reg_64bit_22th_lo,
        // input wire [31:0]                       i_reg_64bit_23th_hi,
        // input wire [31:0]                       i_reg_64bit_23th_lo,
        // input wire [31:0]                       i_reg_64bit_24th_hi,
        // input wire [31:0]                       i_reg_64bit_24th_lo,
        // input wire [31:0]                       i_reg_64bit_25th_hi,
        // input wire [31:0]                       i_reg_64bit_25th_lo,
        // input wire [31:0]                       i_reg_64bit_26th_hi,
        // input wire [31:0]                       i_reg_64bit_26th_lo,
        // input wire [31:0]                       i_reg_64bit_27th_hi,
        // input wire [31:0]                       i_reg_64bit_27th_lo,
        // input wire [31:0]                       i_reg_64bit_28th_hi,
        // input wire [31:0]                       i_reg_64bit_28th_lo,
        // input wire [31:0]                       i_reg_64bit_29th_hi,
        // input wire [31:0]                       i_reg_64bit_29th_lo,
        // input wire [31:0]                       i_reg_64bit_30th_hi,
        // input wire [31:0]                       i_reg_64bit_30th_lo,
        // input wire [31:0]                       i_reg_64bit_31th_hi,
        // input wire [31:0]                       i_reg_64bit_31th_lo,
        // input wire [31:0]                       i_reg_64bit_32th_hi,
        // input wire [31:0]                       i_reg_64bit_32th_lo,
        // input wire [31:0]                       i_reg_64bit_33th_hi,
        // input wire [31:0]                       i_reg_64bit_33th_lo,
        // input wire [31:0]                       i_reg_64bit_34th_hi,
        // input wire [31:0]                       i_reg_64bit_34th_lo,
        // input wire [31:0]                       i_reg_64bit_35th_hi,
        // input wire [31:0]                       i_reg_64bit_35th_lo,
        // input wire [31:0]                       i_reg_64bit_36th_hi,
        // input wire [31:0]                       i_reg_64bit_36th_lo,
        // input wire [31:0]                       i_reg_64bit_37th_hi,
        // input wire [31:0]                       i_reg_64bit_37th_lo,
        // input wire [31:0]                       i_reg_64bit_38th_hi,
        // input wire [31:0]                       i_reg_64bit_38th_lo,
        // input wire [31:0]                       i_reg_64bit_39th_hi,
        // input wire [31:0]                       i_reg_64bit_39th_lo,
        // input wire [31:0]                       i_reg_64bit_40th_hi,
        // input wire [31:0]                       i_reg_64bit_40th_lo,
        // input wire [31:0]                       i_reg_64bit_41th_hi,
        // input wire [31:0]                       i_reg_64bit_41th_lo,
        // input wire [31:0]                       i_reg_64bit_42th_hi,
        // input wire [31:0]                       i_reg_64bit_42th_lo,
        // input wire [31:0]                       i_reg_64bit_43th_hi,
        // input wire [31:0]                       i_reg_64bit_43th_lo,
        // input wire [31:0]                       i_reg_64bit_44th_hi,
        // input wire [31:0]                       i_reg_64bit_44th_lo,
        // input wire [31:0]                       i_reg_64bit_45th_hi,
        // input wire [31:0]                       i_reg_64bit_45th_lo,
        // input wire [31:0]                       i_reg_64bit_46th_hi,
        // input wire [31:0]                       i_reg_64bit_46th_lo,
        // input wire [31:0]                       i_reg_64bit_47th_hi,
        // input wire [31:0]                       i_reg_64bit_47th_lo,
        // input wire [31:0]                       i_reg_64bit_48th_hi,
        // input wire [31:0]                       i_reg_64bit_48th_lo,
        // input wire [31:0]                       i_reg_64bit_49th_hi,
        // input wire [31:0]                       i_reg_64bit_49th_lo,
        // input wire [31:0]                       i_reg_64bit_50th_hi,
        // input wire [31:0]                       i_reg_64bit_50th_lo,
        // input wire [31:0]                       i_reg_64bit_51th_hi,
        // input wire [31:0]                       i_reg_64bit_51th_lo,
        // input wire [31:0]                       i_reg_64bit_52th_hi,
        // input wire [31:0]                       i_reg_64bit_52th_lo,
        // input wire [31:0]                       i_reg_64bit_53th_hi,
        // input wire [31:0]                       i_reg_64bit_53th_lo,
        // input wire [31:0]                       i_reg_64bit_54th_hi,
        // input wire [31:0]                       i_reg_64bit_54th_lo,
        // input wire [31:0]                       i_reg_64bit_55th_hi,
        // input wire [31:0]                       i_reg_64bit_55th_lo,
        // input wire [31:0]                       i_reg_64bit_56th_hi,
        // input wire [31:0]                       i_reg_64bit_56th_lo,
        // input wire [31:0]                       i_reg_64bit_57th_hi,
        // input wire [31:0]                       i_reg_64bit_57th_lo,
        // input wire [31:0]                       i_reg_64bit_58th_hi,
        // input wire [31:0]                       i_reg_64bit_58th_lo,
        // input wire [31:0]                       i_reg_64bit_59th_hi,
        // input wire [31:0]                       i_reg_64bit_59th_lo,
        // input wire [31:0]                       i_reg_64bit_60th_hi,
        // input wire [31:0]                       i_reg_64bit_60th_lo,
        // input wire [31:0]                       i_reg_64bit_61th_hi,
        // input wire [31:0]                       i_reg_64bit_61th_lo,
        // input wire [31:0]                       i_reg_64bit_62th_hi,
        // input wire [31:0]                       i_reg_64bit_62th_lo,
        // input wire [31:0]                       i_reg_64bit_63th_hi,
        // input wire [31:0]                       i_reg_64bit_63th_lo,
        // input wire [31:0]                       i_reg_64bit_64th_hi,
        // input wire [31:0]                       i_reg_64bit_64th_lo,
        // input wire [31:0]                       i_reg_64bit_65th_hi,
        // input wire [31:0]                       i_reg_64bit_65th_lo,
        // input wire [31:0]                       i_reg_64bit_66th_hi,
        // input wire [31:0]                       i_reg_64bit_66th_lo,
        // input wire [31:0]                       i_reg_64bit_67th_hi,
        // input wire [31:0]                       i_reg_64bit_67th_lo,
        // input wire [31:0]                       i_reg_64bit_68th_hi,
        // input wire [31:0]                       i_reg_64bit_68th_lo,
        // input wire [31:0]                       i_reg_64bit_69th_hi,
        // input wire [31:0]                       i_reg_64bit_69th_lo,
        // input wire [31:0]                       i_reg_64bit_70th_hi,
        // input wire [31:0]                       i_reg_64bit_70th_lo,
        // input wire [31:0]                       i_reg_64bit_71th_hi,
        // input wire [31:0]                       i_reg_64bit_71th_lo,
        // input wire [31:0]                       i_reg_64bit_72th_hi,
        // input wire [31:0]                       i_reg_64bit_72th_lo,
        // input wire [31:0]                       i_reg_64bit_73th_hi,
        // input wire [31:0]                       i_reg_64bit_73th_lo,
        // input wire [31:0]                       i_reg_64bit_74th_hi,
        // input wire [31:0]                       i_reg_64bit_74th_lo,
        // input wire [31:0]                       i_reg_64bit_75th_hi,
        // input wire [31:0]                       i_reg_64bit_75th_lo,
        // input wire [31:0]                       i_reg_64bit_76th_hi,
        // input wire [31:0]                       i_reg_64bit_76th_lo,
        // input wire [31:0]                       i_reg_64bit_77th_hi,
        // input wire [31:0]                       i_reg_64bit_77th_lo,
        // input wire [31:0]                       i_reg_64bit_78th_hi,
        // input wire [31:0]                       i_reg_64bit_78th_lo,
        // input wire [31:0]                       i_reg_64bit_79th_hi,
        // input wire [31:0]                       i_reg_64bit_79th_lo,
        // input wire [31:0]                       i_reg_64bit_80th_hi,
        // input wire [31:0]                       i_reg_64bit_80th_lo,
        // input wire [31:0]                       i_reg_64bit_81th_hi,
        // input wire [31:0]                       i_reg_64bit_81th_lo,
        // input wire [31:0]                       i_reg_64bit_82th_hi,
        // input wire [31:0]                       i_reg_64bit_82th_lo,
        // input wire [31:0]                       i_reg_64bit_83th_hi,
        // input wire [31:0]                       i_reg_64bit_83th_lo,
        // input wire [31:0]                       i_reg_64bit_84th_hi,
        // input wire [31:0]                       i_reg_64bit_84th_lo,
        // input wire [31:0]                       i_reg_64bit_85th_hi,
        // input wire [31:0]                       i_reg_64bit_85th_lo,
        // input wire [31:0]                       i_reg_64bit_86th_hi,
        // input wire [31:0]                       i_reg_64bit_86th_lo,
        // input wire [31:0]                       i_reg_64bit_87th_hi,
        // input wire [31:0]                       i_reg_64bit_87th_lo,
        // input wire [31:0]                       i_reg_64bit_88th_hi,
        // input wire [31:0]                       i_reg_64bit_88th_lo,
        // input wire [31:0]                       i_reg_64bit_89th_hi,
        // input wire [31:0]                       i_reg_64bit_89th_lo,
        // input wire [31:0]                       i_reg_64bit_90th_hi,
        // input wire [31:0]                       i_reg_64bit_90th_lo,
        // input wire [31:0]                       i_reg_64bit_91th_hi,
        // input wire [31:0]                       i_reg_64bit_91th_lo,
        // input wire [31:0]                       i_reg_64bit_92th_hi,
        // input wire [31:0]                       i_reg_64bit_92th_lo,
        // input wire [31:0]                       i_reg_64bit_93th_hi,
        // input wire [31:0]                       i_reg_64bit_93th_lo,
        // input wire [31:0]                       i_reg_64bit_94th_hi,
        // input wire [31:0]                       i_reg_64bit_94th_lo,
        // input wire [31:0]                       i_reg_64bit_95th_hi,
        // input wire [31:0]                       i_reg_64bit_95th_lo,
        // input wire [31:0]                       i_reg_64bit_96th_hi,
        // input wire [31:0]                       i_reg_64bit_96th_lo,
        // input wire [31:0]                       i_reg_64bit_97th_hi,
        // input wire [31:0]                       i_reg_64bit_97th_lo,
        // input wire [31:0]                       i_reg_64bit_98th_hi,
        // input wire [31:0]                       i_reg_64bit_98th_lo,
        // input wire [31:0]                       i_reg_64bit_99th_hi,
        // input wire [31:0]                       i_reg_64bit_99th_lo,
        // input wire [31:0]                       i_reg_64bit_100th_hi,
        // input wire [31:0]                       i_reg_64bit_100th_lo,
        // input wire [31:0]                       i_reg_64bit_101th_hi,
        // input wire [31:0]                       i_reg_64bit_101th_lo,
        // input wire [31:0]                       i_reg_64bit_102th_hi,
        // input wire [31:0]                       i_reg_64bit_102th_lo,
        // input wire [31:0]                       i_reg_64bit_103th_hi,
        // input wire [31:0]                       i_reg_64bit_103th_lo,
        // input wire [31:0]                       i_reg_64bit_104th_hi,
        // input wire [31:0]                       i_reg_64bit_104th_lo,
        // input wire [31:0]                       i_reg_64bit_105th_hi,
        // input wire [31:0]                       i_reg_64bit_105th_lo,
        // input wire [31:0]                       i_reg_64bit_106th_hi,
        // input wire [31:0]                       i_reg_64bit_106th_lo,
        // input wire [31:0]                       i_reg_64bit_107th_hi,
        // input wire [31:0]                       i_reg_64bit_107th_lo,
        // input wire [31:0]                       i_reg_64bit_108th_hi,
        // input wire [31:0]                       i_reg_64bit_108th_lo,
        // input wire [31:0]                       i_reg_64bit_109th_hi,
        // input wire [31:0]                       i_reg_64bit_109th_lo,
        // input wire [31:0]                       i_reg_64bit_110th_hi,
        // input wire [31:0]                       i_reg_64bit_110th_lo,
        // input wire [31:0]                       i_reg_64bit_111th_hi,
        // input wire [31:0]                       i_reg_64bit_111th_lo,
        // input wire [31:0]                       i_reg_64bit_112th_hi,
        // input wire [31:0]                       i_reg_64bit_112th_lo,
        // input wire [31:0]                       i_reg_64bit_113th_hi,
        // input wire [31:0]                       i_reg_64bit_113th_lo,
        // input wire [31:0]                       i_reg_64bit_114th_hi,
        // input wire [31:0]                       i_reg_64bit_114th_lo,
        // input wire [31:0]                       i_reg_64bit_115th_hi,
        // input wire [31:0]                       i_reg_64bit_115th_lo,
        // input wire [31:0]                       i_reg_64bit_116th_hi,
        // input wire [31:0]                       i_reg_64bit_116th_lo,
        // input wire [31:0]                       i_reg_64bit_117th_hi,
        // input wire [31:0]                       i_reg_64bit_117th_lo,
        // input wire [31:0]                       i_reg_64bit_118th_hi,
        // input wire [31:0]                       i_reg_64bit_118th_lo,
        // input wire [31:0]                       i_reg_64bit_119th_hi,
        // input wire [31:0]                       i_reg_64bit_119th_lo,
        // input wire [31:0]                       i_reg_64bit_120th_hi,
        // input wire [31:0]                       i_reg_64bit_120th_lo,
        // input wire [31:0]                       i_reg_64bit_121th_hi,
        // input wire [31:0]                       i_reg_64bit_121th_lo,
        // input wire [31:0]                       i_reg_64bit_122th_hi,
        // input wire [31:0]                       i_reg_64bit_122th_lo,
        // input wire [31:0]                       i_reg_64bit_123th_hi,
        // input wire [31:0]                       i_reg_64bit_123th_lo,
        // input wire [31:0]                       i_reg_64bit_124th_hi,
        // input wire [31:0]                       i_reg_64bit_124th_lo,
        // input wire [31:0]                       i_reg_64bit_125th_hi,
        // input wire [31:0]                       i_reg_64bit_125th_lo,
        // input wire [31:0]                       i_reg_64bit_126th_hi,
        // input wire [31:0]                       i_reg_64bit_126th_lo,
        // input wire [31:0]                       i_reg_64bit_127th_hi,
        // input wire [31:0]                       i_reg_64bit_127th_lo,
        // input wire [31:0]                       i_reg_64bit_128th_hi,        // Match to 'slv_reg254'
        // input wire [31:0]                       i_reg_64bit_128th_lo,        // Match to 'slv_reg255'

        // Add User Output Pins  (# User Guide : Uncomment Pins to Use)
        // output wire [31:0]                      o_reg_64bit_1th_hi,          // Match to 'slv_reg0'
        // output wire [31:0]                      o_reg_64bit_1th_lo,          // Match to 'slv_reg1'
        // output wire [31:0]                      o_reg_64bit_2th_hi,
        // output wire [31:0]                      o_reg_64bit_2th_lo,
        // output wire [31:0]                      o_reg_64bit_3th_hi,
        // output wire [31:0]                      o_reg_64bit_3th_lo,
        // output wire [31:0]                      o_reg_64bit_4th_hi,
        // output wire [31:0]                      o_reg_64bit_4th_lo,
        // output wire [31:0]                      o_reg_64bit_5th_hi,
        // output wire [31:0]                      o_reg_64bit_5th_lo,
        // output wire [31:0]                      o_reg_64bit_6th_hi,
        // output wire [31:0]                      o_reg_64bit_6th_lo,
        // output wire [31:0]                      o_reg_64bit_7th_hi,
        // output wire [31:0]                      o_reg_64bit_7th_lo,
        // output wire [31:0]                      o_reg_64bit_8th_hi,
        // output wire [31:0]                      o_reg_64bit_8th_lo,
        // output wire [31:0]                      o_reg_64bit_9th_hi,
        // output wire [31:0]                      o_reg_64bit_9th_lo,
        // output wire [31:0]                      o_reg_64bit_10th_hi,
        // output wire [31:0]                      o_reg_64bit_10th_lo,
        // output wire [31:0]                      o_reg_64bit_11th_hi,
        // output wire [31:0]                      o_reg_64bit_11th_lo,
        // output wire [31:0]                      o_reg_64bit_12th_hi,
        // output wire [31:0]                      o_reg_64bit_12th_lo,
        // output wire [31:0]                      o_reg_64bit_13th_hi,
        // output wire [31:0]                      o_reg_64bit_13th_lo,
        // output wire [31:0]                      o_reg_64bit_14th_hi,
        // output wire [31:0]                      o_reg_64bit_14th_lo,
        // output wire [31:0]                      o_reg_64bit_15th_hi,
        // output wire [31:0]                      o_reg_64bit_15th_lo,
        // output wire [31:0]                      o_reg_64bit_16th_hi,
        // output wire [31:0]                      o_reg_64bit_16th_lo,
        // output wire [31:0]                      o_reg_64bit_17th_hi,
        // output wire [31:0]                      o_reg_64bit_17th_lo,
        // output wire [31:0]                      o_reg_64bit_18th_hi,
        // output wire [31:0]                      o_reg_64bit_18th_lo,
        // output wire [31:0]                      o_reg_64bit_19th_hi,
        // output wire [31:0]                      o_reg_64bit_19th_lo,
        // output wire [31:0]                      o_reg_64bit_20th_hi,
        // output wire [31:0]                      o_reg_64bit_20th_lo,
        // output wire [31:0]                      o_reg_64bit_21th_hi,
        // output wire [31:0]                      o_reg_64bit_21th_lo,
        // output wire [31:0]                      o_reg_64bit_22th_hi,
        // output wire [31:0]                      o_reg_64bit_22th_lo,
        // output wire [31:0]                      o_reg_64bit_23th_hi,
        // output wire [31:0]                      o_reg_64bit_23th_lo,
        // output wire [31:0]                      o_reg_64bit_24th_hi,
        // output wire [31:0]                      o_reg_64bit_24th_lo,
        // output wire [31:0]                      o_reg_64bit_25th_hi,
        // output wire [31:0]                      o_reg_64bit_25th_lo,
        // output wire [31:0]                      o_reg_64bit_26th_hi,
        // output wire [31:0]                      o_reg_64bit_26th_lo,
        // output wire [31:0]                      o_reg_64bit_27th_hi,
        // output wire [31:0]                      o_reg_64bit_27th_lo,
        // output wire [31:0]                      o_reg_64bit_28th_hi,
        // output wire [31:0]                      o_reg_64bit_28th_lo,
        // output wire [31:0]                      o_reg_64bit_29th_hi,
        // output wire [31:0]                      o_reg_64bit_29th_lo,
        // output wire [31:0]                      o_reg_64bit_30th_hi,
        // output wire [31:0]                      o_reg_64bit_30th_lo,
        // output wire [31:0]                      o_reg_64bit_31th_hi,
        // output wire [31:0]                      o_reg_64bit_31th_lo,
        // output wire [31:0]                      o_reg_64bit_32th_hi,
        // output wire [31:0]                      o_reg_64bit_32th_lo,
        // output wire [31:0]                      o_reg_64bit_33th_hi,
        // output wire [31:0]                      o_reg_64bit_33th_lo,
        // output wire [31:0]                      o_reg_64bit_34th_hi,
        // output wire [31:0]                      o_reg_64bit_34th_lo,
        // output wire [31:0]                      o_reg_64bit_35th_hi,
        // output wire [31:0]                      o_reg_64bit_35th_lo,
        // output wire [31:0]                      o_reg_64bit_36th_hi,
        // output wire [31:0]                      o_reg_64bit_36th_lo,
        // output wire [31:0]                      o_reg_64bit_37th_hi,
        // output wire [31:0]                      o_reg_64bit_37th_lo,
        // output wire [31:0]                      o_reg_64bit_38th_hi,
        // output wire [31:0]                      o_reg_64bit_38th_lo,
        // output wire [31:0]                      o_reg_64bit_39th_hi,
        // output wire [31:0]                      o_reg_64bit_39th_lo,
        // output wire [31:0]                      o_reg_64bit_40th_hi,
        // output wire [31:0]                      o_reg_64bit_40th_lo,
        // output wire [31:0]                      o_reg_64bit_41th_hi,
        // output wire [31:0]                      o_reg_64bit_41th_lo,
        // output wire [31:0]                      o_reg_64bit_42th_hi,
        // output wire [31:0]                      o_reg_64bit_42th_lo,
        // output wire [31:0]                      o_reg_64bit_43th_hi,
        // output wire [31:0]                      o_reg_64bit_43th_lo,
        // output wire [31:0]                      o_reg_64bit_44th_hi,
        // output wire [31:0]                      o_reg_64bit_44th_lo,
        // output wire [31:0]                      o_reg_64bit_45th_hi,
        // output wire [31:0]                      o_reg_64bit_45th_lo,
        // output wire [31:0]                      o_reg_64bit_46th_hi,
        // output wire [31:0]                      o_reg_64bit_46th_lo,
        // output wire [31:0]                      o_reg_64bit_47th_hi,
        // output wire [31:0]                      o_reg_64bit_47th_lo,
        // output wire [31:0]                      o_reg_64bit_48th_hi,
        // output wire [31:0]                      o_reg_64bit_48th_lo,
        // output wire [31:0]                      o_reg_64bit_49th_hi,
        // output wire [31:0]                      o_reg_64bit_49th_lo,
        // output wire [31:0]                      o_reg_64bit_50th_hi,
        // output wire [31:0]                      o_reg_64bit_50th_lo,
        // output wire [31:0]                      o_reg_64bit_51th_hi,
        // output wire [31:0]                      o_reg_64bit_51th_lo,
        // output wire [31:0]                      o_reg_64bit_52th_hi,
        // output wire [31:0]                      o_reg_64bit_52th_lo,
        // output wire [31:0]                      o_reg_64bit_53th_hi,
        // output wire [31:0]                      o_reg_64bit_53th_lo,
        // output wire [31:0]                      o_reg_64bit_54th_hi,
        // output wire [31:0]                      o_reg_64bit_54th_lo,
        // output wire [31:0]                      o_reg_64bit_55th_hi,
        // output wire [31:0]                      o_reg_64bit_55th_lo,
        // output wire [31:0]                      o_reg_64bit_56th_hi,
        // output wire [31:0]                      o_reg_64bit_56th_lo,
        // output wire [31:0]                      o_reg_64bit_57th_hi,
        // output wire [31:0]                      o_reg_64bit_57th_lo,
        // output wire [31:0]                      o_reg_64bit_58th_hi,
        // output wire [31:0]                      o_reg_64bit_58th_lo,
        // output wire [31:0]                      o_reg_64bit_59th_hi,
        // output wire [31:0]                      o_reg_64bit_59th_lo,
        // output wire [31:0]                      o_reg_64bit_60th_hi,
        // output wire [31:0]                      o_reg_64bit_60th_lo,
        // output wire [31:0]                      o_reg_64bit_61th_hi,
        // output wire [31:0]                      o_reg_64bit_61th_lo,
        // output wire [31:0]                      o_reg_64bit_62th_hi,
        // output wire [31:0]                      o_reg_64bit_62th_lo,
        // output wire [31:0]                      o_reg_64bit_63th_hi,
        // output wire [31:0]                      o_reg_64bit_63th_lo,
        // output wire [31:0]                      o_reg_64bit_64th_hi,
        // output wire [31:0]                      o_reg_64bit_64th_lo,
        // output wire [31:0]                      o_reg_64bit_65th_hi,
        // output wire [31:0]                      o_reg_64bit_65th_lo,
        // output wire [31:0]                      o_reg_64bit_66th_hi,
        // output wire [31:0]                      o_reg_64bit_66th_lo,
        // output wire [31:0]                      o_reg_64bit_67th_hi,
        // output wire [31:0]                      o_reg_64bit_67th_lo,
        // output wire [31:0]                      o_reg_64bit_68th_hi,
        // output wire [31:0]                      o_reg_64bit_68th_lo,
        // output wire [31:0]                      o_reg_64bit_69th_hi,
        // output wire [31:0]                      o_reg_64bit_69th_lo,
        // output wire [31:0]                      o_reg_64bit_70th_hi,
        // output wire [31:0]                      o_reg_64bit_70th_lo,
        // output wire [31:0]                      o_reg_64bit_71th_hi,
        // output wire [31:0]                      o_reg_64bit_71th_lo,
        // output wire [31:0]                      o_reg_64bit_72th_hi,
        // output wire [31:0]                      o_reg_64bit_72th_lo,
        // output wire [31:0]                      o_reg_64bit_73th_hi,
        // output wire [31:0]                      o_reg_64bit_73th_lo,
        // output wire [31:0]                      o_reg_64bit_74th_hi,
        // output wire [31:0]                      o_reg_64bit_74th_lo,
        // output wire [31:0]                      o_reg_64bit_75th_hi,
        // output wire [31:0]                      o_reg_64bit_75th_lo,
        // output wire [31:0]                      o_reg_64bit_76th_hi,
        // output wire [31:0]                      o_reg_64bit_76th_lo,
        // output wire [31:0]                      o_reg_64bit_77th_hi,
        // output wire [31:0]                      o_reg_64bit_77th_lo,
        // output wire [31:0]                      o_reg_64bit_78th_hi,
        // output wire [31:0]                      o_reg_64bit_78th_lo,
        // output wire [31:0]                      o_reg_64bit_79th_hi,
        // output wire [31:0]                      o_reg_64bit_79th_lo,
        // output wire [31:0]                      o_reg_64bit_80th_hi,
        // output wire [31:0]                      o_reg_64bit_80th_lo,
        // output wire [31:0]                      o_reg_64bit_81th_hi,
        // output wire [31:0]                      o_reg_64bit_81th_lo,
        // output wire [31:0]                      o_reg_64bit_82th_hi,
        // output wire [31:0]                      o_reg_64bit_82th_lo,
        // output wire [31:0]                      o_reg_64bit_83th_hi,
        // output wire [31:0]                      o_reg_64bit_83th_lo,
        // output wire [31:0]                      o_reg_64bit_84th_hi,
        // output wire [31:0]                      o_reg_64bit_84th_lo,
        // output wire [31:0]                      o_reg_64bit_85th_hi,
        // output wire [31:0]                      o_reg_64bit_85th_lo,
        // output wire [31:0]                      o_reg_64bit_86th_hi,
        // output wire [31:0]                      o_reg_64bit_86th_lo,
        // output wire [31:0]                      o_reg_64bit_87th_hi,
        // output wire [31:0]                      o_reg_64bit_87th_lo,
        // output wire [31:0]                      o_reg_64bit_88th_hi,
        // output wire [31:0]                      o_reg_64bit_88th_lo,
        // output wire [31:0]                      o_reg_64bit_89th_hi,
        // output wire [31:0]                      o_reg_64bit_89th_lo,
        // output wire [31:0]                      o_reg_64bit_90th_hi,
        // output wire [31:0]                      o_reg_64bit_90th_lo,
        // output wire [31:0]                      o_reg_64bit_91th_hi,
        // output wire [31:0]                      o_reg_64bit_91th_lo,
        // output wire [31:0]                      o_reg_64bit_92th_hi,
        // output wire [31:0]                      o_reg_64bit_92th_lo,
        // output wire [31:0]                      o_reg_64bit_93th_hi,
        // output wire [31:0]                      o_reg_64bit_93th_lo,
        // output wire [31:0]                      o_reg_64bit_94th_hi,
        // output wire [31:0]                      o_reg_64bit_94th_lo,
        // output wire [31:0]                      o_reg_64bit_95th_hi,
        // output wire [31:0]                      o_reg_64bit_95th_lo,
        // output wire [31:0]                      o_reg_64bit_96th_hi,
        // output wire [31:0]                      o_reg_64bit_96th_lo,
        // output wire [31:0]                      o_reg_64bit_97th_hi,
        // output wire [31:0]                      o_reg_64bit_97th_lo,
        // output wire [31:0]                      o_reg_64bit_98th_hi,
        // output wire [31:0]                      o_reg_64bit_98th_lo,
        // output wire [31:0]                      o_reg_64bit_99th_hi,
        // output wire [31:0]                      o_reg_64bit_99th_lo,
        // output wire [31:0]                      o_reg_64bit_100th_hi,
        // output wire [31:0]                      o_reg_64bit_100th_lo,
        // output wire [31:0]                      o_reg_64bit_101th_hi,
        // output wire [31:0]                      o_reg_64bit_101th_lo,
        // output wire [31:0]                      o_reg_64bit_102th_hi,
        // output wire [31:0]                      o_reg_64bit_102th_lo,
        // output wire [31:0]                      o_reg_64bit_103th_hi,
        // output wire [31:0]                      o_reg_64bit_103th_lo,
        // output wire [31:0]                      o_reg_64bit_104th_hi,
        // output wire [31:0]                      o_reg_64bit_104th_lo,
        // output wire [31:0]                      o_reg_64bit_105th_hi,
        // output wire [31:0]                      o_reg_64bit_105th_lo,
        // output wire [31:0]                      o_reg_64bit_106th_hi,
        // output wire [31:0]                      o_reg_64bit_106th_lo,
        // output wire [31:0]                      o_reg_64bit_107th_hi,
        // output wire [31:0]                      o_reg_64bit_107th_lo,
        // output wire [31:0]                      o_reg_64bit_108th_hi,
        // output wire [31:0]                      o_reg_64bit_108th_lo,
        // output wire [31:0]                      o_reg_64bit_109th_hi,
        // output wire [31:0]                      o_reg_64bit_109th_lo,
        // output wire [31:0]                      o_reg_64bit_110th_hi,
        // output wire [31:0]                      o_reg_64bit_110th_lo,
        // output wire [31:0]                      o_reg_64bit_111th_hi,
        // output wire [31:0]                      o_reg_64bit_111th_lo,
        // output wire [31:0]                      o_reg_64bit_112th_hi,
        // output wire [31:0]                      o_reg_64bit_112th_lo,
        // output wire [31:0]                      o_reg_64bit_113th_hi,
        // output wire [31:0]                      o_reg_64bit_113th_lo,
        // output wire [31:0]                      o_reg_64bit_114th_hi,
        // output wire [31:0]                      o_reg_64bit_114th_lo,
        // output wire [31:0]                      o_reg_64bit_115th_hi,
        // output wire [31:0]                      o_reg_64bit_115th_lo,
        // output wire [31:0]                      o_reg_64bit_116th_hi,
        // output wire [31:0]                      o_reg_64bit_116th_lo,
        // output wire [31:0]                      o_reg_64bit_117th_hi,
        // output wire [31:0]                      o_reg_64bit_117th_lo,
        // output wire [31:0]                      o_reg_64bit_118th_hi,
        // output wire [31:0]                      o_reg_64bit_118th_lo,
        // output wire [31:0]                      o_reg_64bit_119th_hi,
        // output wire [31:0]                      o_reg_64bit_119th_lo,
        // output wire [31:0]                      o_reg_64bit_120th_hi,
        // output wire [31:0]                      o_reg_64bit_120th_lo,
        // output wire [31:0]                      o_reg_64bit_121th_hi,
        // output wire [31:0]                      o_reg_64bit_121th_lo,
        // output wire [31:0]                      o_reg_64bit_122th_hi,
        // output wire [31:0]                      o_reg_64bit_122th_lo,
        // output wire [31:0]                      o_reg_64bit_123th_hi,
        // output wire [31:0]                      o_reg_64bit_123th_lo,
        // output wire [31:0]                      o_reg_64bit_124th_hi,
        // output wire [31:0]                      o_reg_64bit_124th_lo,
        // output wire [31:0]                      o_reg_64bit_125th_hi,
        // output wire [31:0]                      o_reg_64bit_125th_lo,
        // output wire [31:0]                      o_reg_64bit_126th_hi,
        // output wire [31:0]                      o_reg_64bit_126th_lo,
        // output wire [31:0]                      o_reg_64bit_127th_hi,
        // output wire [31:0]                      o_reg_64bit_127th_lo,
        // output wire [31:0]                      o_reg_64bit_128th_hi,            // Match to 'slv_reg254'
        // output wire [31:0]                      o_reg_64bit_128th_lo,            // Match to 'slv_reg255'
        // End User I/O Pins
	);

// ============================================================================ //
//                                                                              //
//                                 Local Param.                                 //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Local Param. to Define the                                      //
// ==================================================================== //
    localparam integer OPT_MEM_ADDR_BITS = 7;

// ============================================================================ //
//                                                                              //
//                                  Wire & Reg                                  //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Variable used for AXI4-Lite Signal                              //
// ==================================================================== //
	// AXI4-LITE Signals
	reg [C_S_AXI_ADDR_WIDTH-1:0]    axi_awaddr;
	reg  	                        axi_awready;
	reg  	                        axi_wready;
	reg [1:0] 	                    axi_bresp;
	reg  	                        axi_bvalid;
	reg [C_S_AXI_ADDR_WIDTH-1:0] 	axi_araddr;
	reg  	                        axi_arready;
	reg [C_S_AXI_DATA_WIDTH-1:0] 	axi_rdata;
	reg [1:0] 	                    axi_rresp;
	reg  	                        axi_rvalid;

    // I/O Connections Assignments
	assign S_AXI_AWREADY    = axi_awready;
	assign S_AXI_WREADY	    = axi_wready;
	assign S_AXI_BRESP	    = axi_bresp;
	assign S_AXI_BVALID	    = axi_bvalid;
	assign S_AXI_ARREADY	= axi_arready;
	assign S_AXI_RDATA	    = axi_rdata;
	assign S_AXI_RRESP	    = axi_rresp;
	assign S_AXI_RVALID	    = axi_rvalid;

// ==================================================================== //
//  [2] Variable used for Slave Register                                //
// ==================================================================== //
    // Slave Register
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg0;           // Match to 'i/o_reg_64bit_1th_hi' I/O Pin
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg1;           // Match to 'i/o_reg_64bit_1th_lo' I/O Pin
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg2;           // Match to 'i/o_reg_64bit_2th_hi' I/O Pin
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg3;           // Match to 'i/o_reg_64bit_2th_lo' I/O Pin
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg4;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg5;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg6;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg7;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg8;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg9;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg10;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg11;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg12;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg13;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg14;
	reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg15;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg16;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg17;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg18;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg19;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg20;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg21;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg22;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg23;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg24;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg25;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg26;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg27;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg28;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg29;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg30;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg31;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg32;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg33;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg34;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg35;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg36;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg37;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg38;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg39;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg40;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg41;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg42;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg43;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg44;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg45;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg46;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg47;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg48;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg49;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg50;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg51;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg52;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg53;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg54;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg55;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg56;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg57;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg58;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg59;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg60;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg61;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg62;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg63;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg64;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg65;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg66;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg67;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg68;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg69;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg70;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg71;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg72;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg73;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg74;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg75;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg76;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg77;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg78;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg79;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg80;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg81;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg82;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg83;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg84;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg85;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg86;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg87;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg88;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg89;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg90;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg91;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg92;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg93;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg94;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg95;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg96;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg97;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg98;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg99;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg100;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg101;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg102;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg103;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg104;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg105;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg106;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg107;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg108;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg109;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg110;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg111;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg112;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg113;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg114;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg115;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg116;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg117;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg118;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg119;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg120;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg121;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg122;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg123;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg124;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg125;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg126;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg127;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg128;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg129;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg130;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg131;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg132;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg133;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg134;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg135;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg136;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg137;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg138;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg139;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg140;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg141;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg142;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg143;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg144;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg145;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg146;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg147;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg148;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg149;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg150;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg151;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg152;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg153;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg154;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg155;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg156;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg157;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg158;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg159;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg160;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg161;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg162;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg163;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg164;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg165;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg166;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg167;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg168;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg169;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg170;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg171;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg172;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg173;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg174;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg175;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg176;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg177;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg178;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg179;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg180;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg181;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg182;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg183;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg184;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg185;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg186;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg187;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg188;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg189;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg190;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg191;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg192;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg193;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg194;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg195;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg196;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg197;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg198;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg199;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg200;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg201;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg202;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg203;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg204;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg205;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg206;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg207;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg208;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg209;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg210;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg211;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg212;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg213;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg214;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg215;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg216;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg217;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg218;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg219;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg220;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg221;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg222;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg223;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg224;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg225;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg226;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg227;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg228;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg229;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg230;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg231;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg232;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg233;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg234;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg235;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg236;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg237;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg238;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg239;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg240;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg241;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg242;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg243;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg244;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg245;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg246;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg247;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg248;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg249;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg250;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg251;
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg252;         // Match to 'i/o_reg_64bit_127th_hi' I/O Pin
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg253;         // Match to 'i/o_reg_64bit_127th_lo' I/O Pin
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg254;         // Match to 'i/o_reg_64bit_128th_hi' I/O Pin
    reg [C_S_AXI_DATA_WIDTH-1:0]	slv_reg255;         // Match to 'i/o_reg_64bit_128th_lo' I/O Pin
	wire	                        slv_reg_rden;
	wire	                        slv_reg_wren;
	reg [C_S_AXI_DATA_WIDTH-1:0]    reg_data_out;
	integer	                        byte_index;
	reg	                            aw_en;

// ============================================================================ //
//                                                                              //
//                       AXI4-Lite Write Transaction Logic                      //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Seq. Logic for Write Address Channel                            //
// ==================================================================== //
    // 1. AWADDR :
    // Write address is latched when both S_AXI_AWVALID and A_AXI_WVALID are valid.
	always @(posedge S_AXI_ACLK) begin
	    if(S_AXI_ARESETN == 1'b0) begin
	        axi_awaddr <= 0;
	    end 
	    else begin
	        if(~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en) begin
	            axi_awaddr <= S_AXI_AWADDR;     // Write address latching
	        end
	    end 
	end   

    // 2. AWREADY :
    // axi_awready is asserted for one S_AXI_ACLK clock cycle when both S_AXI_AWVALID and S_AXI_WVALID are asserted.
    // axi_awready is de-asserted when reset is low.
	always @(posedge S_AXI_ACLK) begin
	    if(S_AXI_ARESETN == 1'b0) begin
            axi_awready <= 1'b0;
            aw_en <= 1'b1;
        end
	    else begin
	        if(~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en) begin
                axi_awready <= 1'b1;
                aw_en <= 1'b0;
	        end
	        else if(S_AXI_BREADY && axi_bvalid) begin
                aw_en <= 1'b1;
                axi_awready <= 1'b0;
	        end
	        else begin
                axi_awready <= 1'b0;
	        end
	    end 
	end       

// ==================================================================== //
//  [2] Seq. Logic for Write Data Channel                               //
// ==================================================================== //

    // 1. WDATA :
    // The write data is accepted and written to memory mapped registers when axi_awready, S_AXI_AWVALID, axi_wready and S_AXI_WVALID are asserted.
    // Write strobes are used to select byte enables of slave registers while writing.
    // These registers are cleared when reset (active low) is applied.
    // Slave register write enable is asserted when valid address and data are available and the slave is ready to accept the write address and write data.
	assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

	always @(posedge S_AXI_ACLK) begin
        if(S_AXI_ARESETN == 1'b0) begin
            // # User Guide : Comment the Registers which are Read-Only or Un-Used
            slv_reg0 <= 0;
            slv_reg1 <= 0;
            slv_reg2 <= 0;
            slv_reg3 <= 0;
            slv_reg4 <= 0;
            slv_reg5 <= 0;
            slv_reg6 <= 0;
            slv_reg7 <= 0;
            slv_reg8 <= 0;
            slv_reg9 <= 0;
            slv_reg10 <= 0;
            slv_reg11 <= 0;
            slv_reg12 <= 0;
            slv_reg13 <= 0;
            slv_reg14 <= 0;
            slv_reg15 <= 0;
            slv_reg16 <= 0;
            slv_reg17 <= 0;
            slv_reg18 <= 0;
            slv_reg19 <= 0;
            slv_reg20 <= 0;
            slv_reg21 <= 0;
            slv_reg22 <= 0;
            slv_reg23 <= 0;
            slv_reg24 <= 0;
            slv_reg25 <= 0;
            slv_reg26 <= 0;
            slv_reg27 <= 0;
            slv_reg28 <= 0;
            slv_reg29 <= 0;
            slv_reg30 <= 0;
            slv_reg31 <= 0;
            slv_reg32 <= 0;
            slv_reg33 <= 0;
            slv_reg34 <= 0;
            slv_reg35 <= 0;
            slv_reg36 <= 0;
            slv_reg37 <= 0;
            slv_reg38 <= 0;
            slv_reg39 <= 0;
            slv_reg40 <= 0;
            slv_reg41 <= 0;
            slv_reg42 <= 0;
            slv_reg43 <= 0;
            slv_reg44 <= 0;
            slv_reg45 <= 0;
            slv_reg46 <= 0;
            slv_reg47 <= 0;
            slv_reg48 <= 0;
            slv_reg49 <= 0;
            slv_reg50 <= 0;
            slv_reg51 <= 0;
            slv_reg52 <= 0;
            slv_reg53 <= 0;
            slv_reg54 <= 0;
            slv_reg55 <= 0;
            slv_reg56 <= 0;
            slv_reg57 <= 0;
            slv_reg58 <= 0;
            slv_reg59 <= 0;
            slv_reg60 <= 0;
            slv_reg61 <= 0;
            slv_reg62 <= 0;
            slv_reg63 <= 0;
            slv_reg64 <= 0;
            slv_reg65 <= 0;
            slv_reg66 <= 0;
            slv_reg67 <= 0;
            slv_reg68 <= 0;
            slv_reg69 <= 0;
            slv_reg70 <= 0;
            slv_reg71 <= 0;
            slv_reg72 <= 0;
            slv_reg73 <= 0;
            slv_reg74 <= 0;
            slv_reg75 <= 0;
            slv_reg76 <= 0;
            slv_reg77 <= 0;
            slv_reg78 <= 0;
            slv_reg79 <= 0;
            slv_reg80 <= 0;
            slv_reg81 <= 0;
            slv_reg82 <= 0;
            slv_reg83 <= 0;
            slv_reg84 <= 0;
            slv_reg85 <= 0;
            slv_reg86 <= 0;
            slv_reg87 <= 0;
            slv_reg88 <= 0;
            slv_reg89 <= 0;
            slv_reg90 <= 0;
            slv_reg91 <= 0;
            slv_reg92 <= 0;
            slv_reg93 <= 0;
            slv_reg94 <= 0;
            slv_reg95 <= 0;
            slv_reg96 <= 0;
            slv_reg97 <= 0;
            slv_reg98 <= 0;
            slv_reg99 <= 0;
            slv_reg100 <= 0;
            slv_reg101 <= 0;
            slv_reg102 <= 0;
            slv_reg103 <= 0;
            slv_reg104 <= 0;
            slv_reg105 <= 0;
            slv_reg106 <= 0;
            slv_reg107 <= 0;
            slv_reg108 <= 0;
            slv_reg109 <= 0;
            slv_reg110 <= 0;
            slv_reg111 <= 0;
            slv_reg112 <= 0;
            slv_reg113 <= 0;
            slv_reg114 <= 0;
            slv_reg115 <= 0;
            slv_reg116 <= 0;
            slv_reg117 <= 0;
            slv_reg118 <= 0;
            slv_reg119 <= 0;
            slv_reg120 <= 0;
            slv_reg121 <= 0;
            slv_reg122 <= 0;
            slv_reg123 <= 0;
            slv_reg124 <= 0;
            slv_reg125 <= 0;
            slv_reg126 <= 0;
            slv_reg127 <= 0;
            slv_reg128 <= 0;
            slv_reg129 <= 0;
            slv_reg130 <= 0;
            slv_reg131 <= 0;
            slv_reg132 <= 0;
            slv_reg133 <= 0;
            slv_reg134 <= 0;
            slv_reg135 <= 0;
            slv_reg136 <= 0;
            slv_reg137 <= 0;
            slv_reg138 <= 0;
            slv_reg139 <= 0;
            slv_reg140 <= 0;
            slv_reg141 <= 0;
            slv_reg142 <= 0;
            slv_reg143 <= 0;
            slv_reg144 <= 0;
            slv_reg145 <= 0;
            slv_reg146 <= 0;
            slv_reg147 <= 0;
            slv_reg148 <= 0;
            slv_reg149 <= 0;
            slv_reg150 <= 0;
            slv_reg151 <= 0;
            slv_reg152 <= 0;
            slv_reg153 <= 0;
            slv_reg154 <= 0;
            slv_reg155 <= 0;
            slv_reg156 <= 0;
            slv_reg157 <= 0;
            slv_reg158 <= 0;
            slv_reg159 <= 0;
            slv_reg160 <= 0;
            slv_reg161 <= 0;
            slv_reg162 <= 0;
            slv_reg163 <= 0;
            slv_reg164 <= 0;
            slv_reg165 <= 0;
            slv_reg166 <= 0;
            slv_reg167 <= 0;
            slv_reg168 <= 0;
            slv_reg169 <= 0;
            slv_reg170 <= 0;
            slv_reg171 <= 0;
            slv_reg172 <= 0;
            slv_reg173 <= 0;
            slv_reg174 <= 0;
            slv_reg175 <= 0;
            slv_reg176 <= 0;
            slv_reg177 <= 0;
            slv_reg178 <= 0;
            slv_reg179 <= 0;
            slv_reg180 <= 0;
            slv_reg181 <= 0;
            slv_reg182 <= 0;
            slv_reg183 <= 0;
            slv_reg184 <= 0;
            slv_reg185 <= 0;
            slv_reg186 <= 0;
            slv_reg187 <= 0;
            slv_reg188 <= 0;
            slv_reg189 <= 0;
            slv_reg190 <= 0;
            slv_reg191 <= 0;
            slv_reg192 <= 0;
            slv_reg193 <= 0;
            slv_reg194 <= 0;
            slv_reg195 <= 0;
            slv_reg196 <= 0;
            slv_reg197 <= 0;
            slv_reg198 <= 0;
            slv_reg199 <= 0;
            slv_reg200 <= 0;
            slv_reg201 <= 0;
            slv_reg202 <= 0;
            slv_reg203 <= 0;
            slv_reg204 <= 0;
            slv_reg205 <= 0;
            slv_reg206 <= 0;
            slv_reg207 <= 0;
            slv_reg208 <= 0;
            slv_reg209 <= 0;
            slv_reg210 <= 0;
            slv_reg211 <= 0;
            slv_reg212 <= 0;
            slv_reg213 <= 0;
            slv_reg214 <= 0;
            slv_reg215 <= 0;
            slv_reg216 <= 0;
            slv_reg217 <= 0;
            slv_reg218 <= 0;
            slv_reg219 <= 0;
            slv_reg220 <= 0;
            slv_reg221 <= 0;
            slv_reg222 <= 0;
            slv_reg223 <= 0;
            slv_reg224 <= 0;
            slv_reg225 <= 0;
            slv_reg226 <= 0;
            slv_reg227 <= 0;
            slv_reg228 <= 0;
            slv_reg229 <= 0;
            slv_reg230 <= 0;
            slv_reg231 <= 0;
            slv_reg232 <= 0;
            slv_reg233 <= 0;
            slv_reg234 <= 0;
            slv_reg235 <= 0;
            slv_reg236 <= 0;
            slv_reg237 <= 0;
            slv_reg238 <= 0;
            slv_reg239 <= 0;
            slv_reg240 <= 0;
            slv_reg241 <= 0;
            slv_reg242 <= 0;
            slv_reg243 <= 0;
            slv_reg244 <= 0;
            slv_reg245 <= 0;
            slv_reg246 <= 0;
            slv_reg247 <= 0;
            slv_reg248 <= 0;
            slv_reg249 <= 0;
            slv_reg250 <= 0;
            slv_reg251 <= 0;
            slv_reg252 <= 0;
            slv_reg253 <= 0;
            slv_reg254 <= 0;
            slv_reg255 <= 0;
	    end 
	    else begin
	        if(slv_reg_wren) begin
	            case(axi_awaddr[OPT_MEM_ADDR_BITS+2:2])
                    // # User Guide : Comment the Registers which are Read-Only or Un-Used
                    8'h00:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 0
                                slv_reg0[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h01:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 1
                                slv_reg1[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h02:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 2
                                slv_reg2[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h03:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 3
                                slv_reg3[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h04:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 4
                                slv_reg4[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h05:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 5
                                slv_reg5[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h06:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 6
                                slv_reg6[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h07:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 7
                                slv_reg7[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h08:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 8
                                slv_reg8[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h09:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 9
                                slv_reg9[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 10
                                slv_reg10[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 11
                                slv_reg11[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 12
                                slv_reg12[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 13
                                slv_reg13[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 14
                                slv_reg14[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h0F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 15
                                slv_reg15[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h10:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 16
                                slv_reg16[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h11:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 17
                                slv_reg17[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h12:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 18
                                slv_reg18[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h13:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 19
                                slv_reg19[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h14:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 20
                                slv_reg20[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h15:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 21
                                slv_reg21[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h16:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 22
                                slv_reg22[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h17:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 23
                                slv_reg23[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h18:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 24
                                slv_reg24[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h19:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 25
                                slv_reg25[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 26
                                slv_reg26[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 27
                                slv_reg27[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 28
                                slv_reg28[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 29
                                slv_reg29[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 30
                                slv_reg30[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h1F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 31
                                slv_reg31[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h20:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 32
                                slv_reg32[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h21:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 33
                                slv_reg33[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h22:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 34
                                slv_reg34[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h23:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 35
                                slv_reg35[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h24:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 36
                                slv_reg36[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h25:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 37
                                slv_reg37[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h26:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 38
                                slv_reg38[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h27:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 39
                                slv_reg39[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h28:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 40
                                slv_reg40[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h29:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 41
                                slv_reg41[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 42
                                slv_reg42[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 43
                                slv_reg43[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 44
                                slv_reg44[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 45
                                slv_reg45[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 46
                                slv_reg46[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h2F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 47
                                slv_reg47[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h30:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 48
                                slv_reg48[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h31:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 49
                                slv_reg49[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h32:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 50
                                slv_reg50[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h33:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 51
                                slv_reg51[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h34:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 52
                                slv_reg52[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h35:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 53
                                slv_reg53[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h36:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 54
                                slv_reg54[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h37:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 55
                                slv_reg55[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h38:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 56
                                slv_reg56[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h39:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 57
                                slv_reg57[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 58
                                slv_reg58[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 59
                                slv_reg59[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 60
                                slv_reg60[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 61
                                slv_reg61[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 62
                                slv_reg62[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h3F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 63
                                slv_reg63[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h40:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 64
                                slv_reg64[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h41:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 65
                                slv_reg65[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h42:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 66
                                slv_reg66[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h43:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 67
                                slv_reg67[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h44:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 68
                                slv_reg68[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h45:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 69
                                slv_reg69[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h46:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 70
                                slv_reg70[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h47:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 71
                                slv_reg71[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h48:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 72
                                slv_reg72[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h49:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 73
                                slv_reg73[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 74
                                slv_reg74[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 75
                                slv_reg75[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 76
                                slv_reg76[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 77
                                slv_reg77[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 78
                                slv_reg78[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h4F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 79
                                slv_reg79[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h50:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 80
                                slv_reg80[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h51:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 81
                                slv_reg81[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h52:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 82
                                slv_reg82[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h53:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 83
                                slv_reg83[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h54:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 84
                                slv_reg84[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h55:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 85
                                slv_reg85[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h56:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 86
                                slv_reg86[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h57:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 87
                                slv_reg87[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h58:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 88
                                slv_reg88[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h59:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 89
                                slv_reg89[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 90
                                slv_reg90[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 91
                                slv_reg91[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 92
                                slv_reg92[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 93
                                slv_reg93[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 94
                                slv_reg94[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h5F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 95
                                slv_reg95[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h60:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 96
                                slv_reg96[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h61:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 97
                                slv_reg97[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h62:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 98
                                slv_reg98[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h63:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 99
                                slv_reg99[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h64:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 100
                                slv_reg100[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h65:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 101
                                slv_reg101[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h66:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 102
                                slv_reg102[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h67:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 103
                                slv_reg103[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h68:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 104
                                slv_reg104[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h69:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 105
                                slv_reg105[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 106
                                slv_reg106[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 107
                                slv_reg107[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 108
                                slv_reg108[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 109
                                slv_reg109[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 110
                                slv_reg110[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h6F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 111
                                slv_reg111[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h70:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 112
                                slv_reg112[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h71:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 113
                                slv_reg113[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h72:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 114
                                slv_reg114[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h73:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 115
                                slv_reg115[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h74:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 116
                                slv_reg116[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h75:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 117
                                slv_reg117[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h76:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 118
                                slv_reg118[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h77:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 119
                                slv_reg119[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h78:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 120
                                slv_reg120[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h79:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 121
                                slv_reg121[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 122
                                slv_reg122[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 123
                                slv_reg123[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 124
                                slv_reg124[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 125
                                slv_reg125[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 126
                                slv_reg126[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h7F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 127
                                slv_reg127[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h80:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 128
                                slv_reg128[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h81:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 129
                                slv_reg129[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h82:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 130
                                slv_reg130[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h83:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 131
                                slv_reg131[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h84:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 132
                                slv_reg132[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h85:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 133
                                slv_reg133[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h86:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 134
                                slv_reg134[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h87:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 135
                                slv_reg135[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h88:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 136
                                slv_reg136[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h89:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 137
                                slv_reg137[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 138
                                slv_reg138[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 139
                                slv_reg139[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 140
                                slv_reg140[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 141
                                slv_reg141[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 142
                                slv_reg142[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h8F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 143
                                slv_reg143[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h90:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 144
                                slv_reg144[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h91:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 145
                                slv_reg145[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h92:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 146
                                slv_reg146[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h93:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 147
                                slv_reg147[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h94:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 148
                                slv_reg148[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h95:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 149
                                slv_reg149[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h96:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 150
                                slv_reg150[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h97:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 151
                                slv_reg151[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h98:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 152
                                slv_reg152[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h99:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 153
                                slv_reg153[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9A:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 154
                                slv_reg154[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9B:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 155
                                slv_reg155[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9C:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 156
                                slv_reg156[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9D:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 157
                                slv_reg157[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9E:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 158
                                slv_reg158[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'h9F:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 159
                                slv_reg159[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 160
                                slv_reg160[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 161
                                slv_reg161[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 162
                                slv_reg162[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 163
                                slv_reg163[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 164
                                slv_reg164[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 165
                                slv_reg165[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 166
                                slv_reg166[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 167
                                slv_reg167[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 168
                                slv_reg168[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hA9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 169
                                slv_reg169[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 170
                                slv_reg170[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 171
                                slv_reg171[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 172
                                slv_reg172[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAD:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 173
                                slv_reg173[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 174
                                slv_reg174[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hAF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 175
                                slv_reg175[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 176
                                slv_reg176[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 177
                                slv_reg177[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 178
                                slv_reg178[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 179
                                slv_reg179[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 180
                                slv_reg180[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 181
                                slv_reg181[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 182
                                slv_reg182[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 183
                                slv_reg183[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 184
                                slv_reg184[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hB9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 185
                                slv_reg185[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 186
                                slv_reg186[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 187
                                slv_reg187[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 188
                                slv_reg188[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBD:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 189
                                slv_reg189[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 190
                                slv_reg190[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hBF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 191
                                slv_reg191[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 192
                                slv_reg192[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 193
                                slv_reg193[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 194
                                slv_reg194[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 195
                                slv_reg195[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 196
                                slv_reg196[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 197
                                slv_reg197[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 198
                                slv_reg198[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 199
                                slv_reg199[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 200
                                slv_reg200[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hC9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 201
                                slv_reg201[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 202
                                slv_reg202[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 203
                                slv_reg203[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 204
                                slv_reg204[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCD:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 205
                                slv_reg205[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 206
                                slv_reg206[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hCF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 207
                                slv_reg207[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 208
                                slv_reg208[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 209
                                slv_reg209[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 210
                                slv_reg210[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 211
                                slv_reg211[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 212
                                slv_reg212[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 213
                                slv_reg213[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 214
                                slv_reg214[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 215
                                slv_reg215[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 216
                                slv_reg216[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hD9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 217
                                slv_reg217[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 218
                                slv_reg218[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 219
                                slv_reg219[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 220
                                slv_reg220[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDD:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 221
                                slv_reg221[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 222
                                slv_reg222[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hDF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 223
                                slv_reg223[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 224
                                slv_reg224[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 225
                                slv_reg225[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 226
                                slv_reg226[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 227
                                slv_reg227[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 228
                                slv_reg228[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 229
                                slv_reg229[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 230
                                slv_reg230[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 231
                                slv_reg231[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 232
                                slv_reg232[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hE9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 233
                                slv_reg233[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hEA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 234
                                slv_reg234[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hEB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 235
                                slv_reg235[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hEC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 236
                                slv_reg236[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hED:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 237
                                slv_reg237[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hEE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 238
                                slv_reg238[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hEF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 239
                                slv_reg239[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF0:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 240
                                slv_reg240[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF1:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 241
                                slv_reg241[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF2:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 242
                                slv_reg242[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF3:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 243
                                slv_reg243[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF4:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 244
                                slv_reg244[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF5:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 245
                                slv_reg245[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF6:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 246
                                slv_reg246[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF7:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 247
                                slv_reg247[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF8:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 248
                                slv_reg248[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hF9:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 249
                                slv_reg249[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFA:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 250
                                slv_reg250[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFB:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 251
                                slv_reg251[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFC:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 252
                                slv_reg252[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFD:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 253
                                slv_reg253[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFE:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 254
                                slv_reg254[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    8'hFF:
                        for(byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1)
                            if(S_AXI_WSTRB[byte_index] == 1) begin
                                // Respective byte enables are asserted as per write strobes 
                                // Slave register 255
                                slv_reg255[(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
                            end  
                    default :   begin
                                    // # User Guide : Comment the Registers which are Read-Only or Un-Used
                                    slv_reg0 <= slv_reg0;
                                    slv_reg1 <= slv_reg1;
                                    slv_reg2 <= slv_reg2;
                                    slv_reg3 <= slv_reg3;
                                    slv_reg4 <= slv_reg4;
                                    slv_reg5 <= slv_reg5;
                                    slv_reg6 <= slv_reg6;           
                                    slv_reg7 <= slv_reg7;
                                    slv_reg8 <= slv_reg8;
                                    slv_reg9 <= slv_reg9;
                                    slv_reg10 <= slv_reg10;
                                    slv_reg11 <= slv_reg11;
                                    slv_reg12 <= slv_reg12;
                                    slv_reg13 <= slv_reg13;
                                    slv_reg14 <= slv_reg14;
                                    slv_reg15 <= slv_reg15;
                                    slv_reg16 <= slv_reg16;
                                    slv_reg17 <= slv_reg17;
                                    slv_reg18 <= slv_reg18;
                                    slv_reg19 <= slv_reg19;
                                    slv_reg20 <= slv_reg20;
                                    slv_reg21 <= slv_reg21;
                                    slv_reg22 <= slv_reg22;
                                    slv_reg23 <= slv_reg23;
                                    slv_reg24 <= slv_reg24;
                                    slv_reg25 <= slv_reg25;
                                    slv_reg26 <= slv_reg26;
                                    slv_reg27 <= slv_reg27;
                                    slv_reg28 <= slv_reg28;
                                    slv_reg29 <= slv_reg29;
                                    slv_reg30 <= slv_reg30;
                                    slv_reg31 <= slv_reg31;
                                    slv_reg32 <= slv_reg32;
                                    slv_reg33 <= slv_reg33;
                                    slv_reg34 <= slv_reg34;
                                    slv_reg35 <= slv_reg35;
                                    slv_reg36 <= slv_reg36;
                                    slv_reg37 <= slv_reg37;
                                    slv_reg38 <= slv_reg38;
                                    slv_reg39 <= slv_reg39;
                                    slv_reg40 <= slv_reg40;
                                    slv_reg41 <= slv_reg41;
                                    slv_reg42 <= slv_reg42;
                                    slv_reg43 <= slv_reg43;
                                    slv_reg44 <= slv_reg44;
                                    slv_reg45 <= slv_reg45;
                                    slv_reg46 <= slv_reg46;
                                    slv_reg47 <= slv_reg47;
                                    slv_reg48 <= slv_reg48;
                                    slv_reg49 <= slv_reg49;
                                    slv_reg50 <= slv_reg50;
                                    slv_reg51 <= slv_reg51;
                                    slv_reg52 <= slv_reg52;
                                    slv_reg53 <= slv_reg53;
                                    slv_reg54 <= slv_reg54;
                                    slv_reg55 <= slv_reg55;
                                    slv_reg56 <= slv_reg56;
                                    slv_reg57 <= slv_reg57;
                                    slv_reg58 <= slv_reg58;
                                    slv_reg59 <= slv_reg59;
                                    slv_reg60 <= slv_reg60;
                                    slv_reg61 <= slv_reg61;
                                    slv_reg62 <= slv_reg62;
                                    slv_reg63 <= slv_reg63;
                                    slv_reg64 <= slv_reg64;
                                    slv_reg65 <= slv_reg65;
                                    slv_reg66 <= slv_reg66;
                                    slv_reg67 <= slv_reg67;
                                    slv_reg68 <= slv_reg68;
                                    slv_reg69 <= slv_reg69;
                                    slv_reg70 <= slv_reg70;
                                    slv_reg71 <= slv_reg71;
                                    slv_reg72 <= slv_reg72;
                                    slv_reg73 <= slv_reg73;
                                    slv_reg74 <= slv_reg74;
                                    slv_reg75 <= slv_reg75;
                                    slv_reg76 <= slv_reg76;
                                    slv_reg77 <= slv_reg77;
                                    slv_reg78 <= slv_reg78;
                                    slv_reg79 <= slv_reg79;
                                    slv_reg80 <= slv_reg80;
                                    slv_reg81 <= slv_reg81;
                                    slv_reg82 <= slv_reg82;
                                    slv_reg83 <= slv_reg83;
                                    slv_reg84 <= slv_reg84;
                                    slv_reg85 <= slv_reg85;
                                    slv_reg86 <= slv_reg86;
                                    slv_reg87 <= slv_reg87;
                                    slv_reg88 <= slv_reg88;
                                    slv_reg89 <= slv_reg89;
                                    slv_reg90 <= slv_reg90;
                                    slv_reg91 <= slv_reg91;
                                    slv_reg92 <= slv_reg92;
                                    slv_reg93 <= slv_reg93;
                                    slv_reg94 <= slv_reg94;
                                    slv_reg95 <= slv_reg95;
                                    slv_reg96 <= slv_reg96;
                                    slv_reg97 <= slv_reg97;
                                    slv_reg98 <= slv_reg98;
                                    slv_reg99 <= slv_reg99;
                                    slv_reg100 <= slv_reg100;
                                    slv_reg101 <= slv_reg101;
                                    slv_reg102 <= slv_reg102;
                                    slv_reg103 <= slv_reg103;
                                    slv_reg104 <= slv_reg104;
                                    slv_reg105 <= slv_reg105;
                                    slv_reg106 <= slv_reg106;
                                    slv_reg107 <= slv_reg107;
                                    slv_reg108 <= slv_reg108;
                                    slv_reg109 <= slv_reg109;
                                    slv_reg110 <= slv_reg110;
                                    slv_reg111 <= slv_reg111;
                                    slv_reg112 <= slv_reg112;
                                    slv_reg113 <= slv_reg113;
                                    slv_reg114 <= slv_reg114;
                                    slv_reg115 <= slv_reg115;
                                    slv_reg116 <= slv_reg116;
                                    slv_reg117 <= slv_reg117;
                                    slv_reg118 <= slv_reg118;
                                    slv_reg119 <= slv_reg119;
                                    slv_reg120 <= slv_reg120;
                                    slv_reg121 <= slv_reg121;
                                    slv_reg122 <= slv_reg122;
                                    slv_reg123 <= slv_reg123;
                                    slv_reg124 <= slv_reg124;
                                    slv_reg125 <= slv_reg125;
                                    slv_reg126 <= slv_reg126;
                                    slv_reg127 <= slv_reg127;
                                    slv_reg128 <= slv_reg128;
                                    slv_reg129 <= slv_reg129;
                                    slv_reg130 <= slv_reg130;
                                    slv_reg131 <= slv_reg131;
                                    slv_reg132 <= slv_reg132;
                                    slv_reg133 <= slv_reg133;
                                    slv_reg134 <= slv_reg134;
                                    slv_reg135 <= slv_reg135;
                                    slv_reg136 <= slv_reg136;
                                    slv_reg137 <= slv_reg137;
                                    slv_reg138 <= slv_reg138;
                                    slv_reg139 <= slv_reg139;
                                    slv_reg140 <= slv_reg140;
                                    slv_reg141 <= slv_reg141;
                                    slv_reg142 <= slv_reg142;
                                    slv_reg143 <= slv_reg143;
                                    slv_reg144 <= slv_reg144;
                                    slv_reg145 <= slv_reg145;
                                    slv_reg146 <= slv_reg146;
                                    slv_reg147 <= slv_reg147;
                                    slv_reg148 <= slv_reg148;
                                    slv_reg149 <= slv_reg149;
                                    slv_reg150 <= slv_reg150;
                                    slv_reg151 <= slv_reg151;
                                    slv_reg152 <= slv_reg152;
                                    slv_reg153 <= slv_reg153;
                                    slv_reg154 <= slv_reg154;
                                    slv_reg155 <= slv_reg155;
                                    slv_reg156 <= slv_reg156;
                                    slv_reg157 <= slv_reg157;
                                    slv_reg158 <= slv_reg158;
                                    slv_reg159 <= slv_reg159;
                                    slv_reg160 <= slv_reg160;
                                    slv_reg161 <= slv_reg161;
                                    slv_reg162 <= slv_reg162;
                                    slv_reg163 <= slv_reg163;
                                    slv_reg164 <= slv_reg164;
                                    slv_reg165 <= slv_reg165;
                                    slv_reg166 <= slv_reg166;
                                    slv_reg167 <= slv_reg167;
                                    slv_reg168 <= slv_reg168;
                                    slv_reg169 <= slv_reg169;
                                    slv_reg170 <= slv_reg170;
                                    slv_reg171 <= slv_reg171;
                                    slv_reg172 <= slv_reg172;
                                    slv_reg173 <= slv_reg173;
                                    slv_reg174 <= slv_reg174;
                                    slv_reg175 <= slv_reg175;
                                    slv_reg176 <= slv_reg176;
                                    slv_reg177 <= slv_reg177;
                                    slv_reg178 <= slv_reg178;
                                    slv_reg179 <= slv_reg179;
                                    slv_reg180 <= slv_reg180;
                                    slv_reg181 <= slv_reg181;
                                    slv_reg182 <= slv_reg182;
                                    slv_reg183 <= slv_reg183;
                                    slv_reg184 <= slv_reg184;
                                    slv_reg185 <= slv_reg185;
                                    slv_reg186 <= slv_reg186;
                                    slv_reg187 <= slv_reg187;
                                    slv_reg188 <= slv_reg188;
                                    slv_reg189 <= slv_reg189;
                                    slv_reg190 <= slv_reg190;
                                    slv_reg191 <= slv_reg191;
                                    slv_reg192 <= slv_reg192;
                                    slv_reg193 <= slv_reg193;
                                    slv_reg194 <= slv_reg194;
                                    slv_reg195 <= slv_reg195;
                                    slv_reg196 <= slv_reg196;
                                    slv_reg197 <= slv_reg197;
                                    slv_reg198 <= slv_reg198;
                                    slv_reg199 <= slv_reg199;
                                    slv_reg200 <= slv_reg200;
                                    slv_reg201 <= slv_reg201;
                                    slv_reg202 <= slv_reg202;
                                    slv_reg203 <= slv_reg203;
                                    slv_reg204 <= slv_reg204;
                                    slv_reg205 <= slv_reg205;
                                    slv_reg206 <= slv_reg206;
                                    slv_reg207 <= slv_reg207;
                                    slv_reg208 <= slv_reg208;
                                    slv_reg209 <= slv_reg209;
                                    slv_reg210 <= slv_reg210;
                                    slv_reg211 <= slv_reg211;
                                    slv_reg212 <= slv_reg212;
                                    slv_reg213 <= slv_reg213;
                                    slv_reg214 <= slv_reg214;
                                    slv_reg215 <= slv_reg215;
                                    slv_reg216 <= slv_reg216;
                                    slv_reg217 <= slv_reg217;
                                    slv_reg218 <= slv_reg218;
                                    slv_reg219 <= slv_reg219;
                                    slv_reg220 <= slv_reg220;
                                    slv_reg221 <= slv_reg221;
                                    slv_reg222 <= slv_reg222;
                                    slv_reg223 <= slv_reg223;
                                    slv_reg224 <= slv_reg224;
                                    slv_reg225 <= slv_reg225;
                                    slv_reg226 <= slv_reg226;
                                    slv_reg227 <= slv_reg227;
                                    slv_reg228 <= slv_reg228;
                                    slv_reg229 <= slv_reg229;
                                    slv_reg230 <= slv_reg230;
                                    slv_reg231 <= slv_reg231;
                                    slv_reg232 <= slv_reg232;
                                    slv_reg233 <= slv_reg233;
                                    slv_reg234 <= slv_reg234;
                                    slv_reg235 <= slv_reg235;
                                    slv_reg236 <= slv_reg236;
                                    slv_reg237 <= slv_reg237;
                                    slv_reg238 <= slv_reg238;
                                    slv_reg239 <= slv_reg239;
                                    slv_reg240 <= slv_reg240;
                                    slv_reg241 <= slv_reg241;
                                    slv_reg242 <= slv_reg242;
                                    slv_reg243 <= slv_reg243;
                                    slv_reg244 <= slv_reg244;
                                    slv_reg245 <= slv_reg245;
                                    slv_reg246 <= slv_reg246;
                                    slv_reg247 <= slv_reg247;
                                    slv_reg248 <= slv_reg248;
                                    slv_reg249 <= slv_reg249;
                                    slv_reg250 <= slv_reg250;
                                    slv_reg251 <= slv_reg251;
                                    slv_reg252 <= slv_reg252;
                                    slv_reg253 <= slv_reg253;
                                    slv_reg254 <= slv_reg254;
                                    slv_reg255 <= slv_reg255;
                                end
                endcase
	        end
	    end
	end  


    // 2. WREADY :
    // axi_wready is asserted for one S_AXI_ACLK clock cycle when both S_AXI_AWVALID and S_AXI_WVALID are asserted.
	// axi_wready is de-asserted when reset is low.
	always @(posedge S_AXI_ACLK) begin
	    if(S_AXI_ARESETN == 1'b0) begin
	        axi_wready <= 1'b0;
	    end 
	    else begin	        
	        if(~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en) begin
                axi_wready <= 1'b1;
	        end
	        else begin
	            axi_wready <= 1'b0;
	        end
	    end 
	end       

// ==================================================================== //
//  [3] Seq. Logic for Write Response Channel                           //
// ==================================================================== //

    // 1. BVALID & BRESP :
    // The write response and response valid signals are asserted by the slave when axi_awready, S_AXI_AWVALID, axi_wready and S_AXI_WVALID are asserted.
    // This marks the acceptance of address and indicates the status of write transaction.
	always @(posedge S_AXI_ACLK) begin
	    if(S_AXI_ARESETN == 1'b0) begin
            axi_bvalid  <= 0;
            axi_bresp   <= 2'b0;
	    end 
	    else begin
	        if(axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID) begin
                // indicates a valid write response is available
                axi_bvalid <= 1'b1;
                axi_bresp  <= 2'b0; // 'OKAY' response 
	        end
	        else begin
	            if(S_AXI_BREADY && axi_bvalid) begin
                    //check if bready is asserted while bvalid is high) 
                    //(there is a possibility that bready is always asserted high)   
                    axi_bvalid <= 1'b0; 
	            end  
	        end
	    end
	end   

// ============================================================================ //
//                                                                              //
//                       AXI4-Lite Read Transaction Logic                       //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Seq. Logic for Read Address Channel                             //
// ==================================================================== //

    // 1. ARADDR & ARREADY :
    // The read address is also latched when S_AXI_ARVALID is asserted.
    // axi_araddr is reset to zero on reset assertion.
    // axi_arready is asserted for one S_AXI_ACLK clock cycle when S_AXI_ARVALID is asserted.
    // axi_arready is de-asserted when reset (active low) is asserted.
	always @(posedge S_AXI_ACLK) begin
	    if(S_AXI_ARESETN == 1'b0) begin
	        axi_arready <= 1'b0;
	        axi_araddr  <= 32'b0;
	    end 
	    else begin
	        if(~axi_arready && S_AXI_ARVALID) begin
	            // indicates that the slave has acceped the valid read address
	            axi_arready <= 1'b1;
	            // Read address latching
	            axi_araddr  <= S_AXI_ARADDR;
	        end
	        else begin
	            axi_arready <= 1'b0;
	        end
	    end 
	end       

// ==================================================================== //
//  [2] Seq. Logic for Read Data Channel                                //
// ==================================================================== //

    // 1. RDATA :
    // Slave register read enable is asserted when valid address is available and the slave is ready to accept the read address.
	assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;

	always @(*) begin
        // Address decoding for reading registers
        case(axi_araddr[OPT_MEM_ADDR_BITS+2:2])
            8'h00   : reg_data_out <= slv_reg0;
	        8'h01   : reg_data_out <= slv_reg1;
	        8'h02   : reg_data_out <= slv_reg2;
	        8'h03   : reg_data_out <= slv_reg3;
	        8'h04   : reg_data_out <= slv_reg4;
	        8'h05   : reg_data_out <= slv_reg5;
	        8'h06   : reg_data_out <= slv_reg6;
	        8'h07   : reg_data_out <= slv_reg7;
	        8'h08   : reg_data_out <= slv_reg8;
	        8'h09   : reg_data_out <= slv_reg9;
	        8'h0A   : reg_data_out <= slv_reg10;
	        8'h0B   : reg_data_out <= slv_reg11;
	        8'h0C   : reg_data_out <= slv_reg12;
	        8'h0D   : reg_data_out <= slv_reg13;
	        8'h0E   : reg_data_out <= slv_reg14;
	        8'h0F   : reg_data_out <= slv_reg15;
	        8'h10   : reg_data_out <= slv_reg16;
	        8'h11   : reg_data_out <= slv_reg17;
	        8'h12   : reg_data_out <= slv_reg18;
	        8'h13   : reg_data_out <= slv_reg19;
	        8'h14   : reg_data_out <= slv_reg20;
	        8'h15   : reg_data_out <= slv_reg21;
	        8'h16   : reg_data_out <= slv_reg22;
	        8'h17   : reg_data_out <= slv_reg23;
	        8'h18   : reg_data_out <= slv_reg24;
	        8'h19   : reg_data_out <= slv_reg25;
	        8'h1A   : reg_data_out <= slv_reg26;
	        8'h1B   : reg_data_out <= slv_reg27;
	        8'h1C   : reg_data_out <= slv_reg28;
	        8'h1D   : reg_data_out <= slv_reg29;
	        8'h1E   : reg_data_out <= slv_reg30;
	        8'h1F   : reg_data_out <= slv_reg31;
	        8'h20   : reg_data_out <= slv_reg32;
	        8'h21   : reg_data_out <= slv_reg33;
	        8'h22   : reg_data_out <= slv_reg34;
	        8'h23   : reg_data_out <= slv_reg35;
	        8'h24   : reg_data_out <= slv_reg36;
	        8'h25   : reg_data_out <= slv_reg37;
	        8'h26   : reg_data_out <= slv_reg38;
	        8'h27   : reg_data_out <= slv_reg39;
	        8'h28   : reg_data_out <= slv_reg40;
	        8'h29   : reg_data_out <= slv_reg41;
	        8'h2A   : reg_data_out <= slv_reg42;
	        8'h2B   : reg_data_out <= slv_reg43;
	        8'h2C   : reg_data_out <= slv_reg44;
	        8'h2D   : reg_data_out <= slv_reg45;
	        8'h2E   : reg_data_out <= slv_reg46;
	        8'h2F   : reg_data_out <= slv_reg47;
	        8'h30   : reg_data_out <= slv_reg48;
	        8'h31   : reg_data_out <= slv_reg49;
	        8'h32   : reg_data_out <= slv_reg50;
	        8'h33   : reg_data_out <= slv_reg51;
	        8'h34   : reg_data_out <= slv_reg52;
	        8'h35   : reg_data_out <= slv_reg53;
	        8'h36   : reg_data_out <= slv_reg54;
	        8'h37   : reg_data_out <= slv_reg55;
	        8'h38   : reg_data_out <= slv_reg56;
	        8'h39   : reg_data_out <= slv_reg57;
	        8'h3A   : reg_data_out <= slv_reg58;
	        8'h3B   : reg_data_out <= slv_reg59;
	        8'h3C   : reg_data_out <= slv_reg60;
	        8'h3D   : reg_data_out <= slv_reg61;
	        8'h3E   : reg_data_out <= slv_reg62;
	        8'h3F   : reg_data_out <= slv_reg63;
	        8'h40   : reg_data_out <= slv_reg64;
	        8'h41   : reg_data_out <= slv_reg65;
	        8'h42   : reg_data_out <= slv_reg66;
	        8'h43   : reg_data_out <= slv_reg67;
	        8'h44   : reg_data_out <= slv_reg68;
	        8'h45   : reg_data_out <= slv_reg69;
	        8'h46   : reg_data_out <= slv_reg70;
	        8'h47   : reg_data_out <= slv_reg71;
	        8'h48   : reg_data_out <= slv_reg72;
	        8'h49   : reg_data_out <= slv_reg73;
	        8'h4A   : reg_data_out <= slv_reg74;
	        8'h4B   : reg_data_out <= slv_reg75;
	        8'h4C   : reg_data_out <= slv_reg76;
	        8'h4D   : reg_data_out <= slv_reg77;
	        8'h4E   : reg_data_out <= slv_reg78;
	        8'h4F   : reg_data_out <= slv_reg79;
	        8'h50   : reg_data_out <= slv_reg80;
	        8'h51   : reg_data_out <= slv_reg81;
	        8'h52   : reg_data_out <= slv_reg82;
	        8'h53   : reg_data_out <= slv_reg83;
	        8'h54   : reg_data_out <= slv_reg84;
	        8'h55   : reg_data_out <= slv_reg85;
	        8'h56   : reg_data_out <= slv_reg86;
	        8'h57   : reg_data_out <= slv_reg87;
	        8'h58   : reg_data_out <= slv_reg88;
	        8'h59   : reg_data_out <= slv_reg89;
	        8'h5A   : reg_data_out <= slv_reg90;
	        8'h5B   : reg_data_out <= slv_reg91;
	        8'h5C   : reg_data_out <= slv_reg92;
	        8'h5D   : reg_data_out <= slv_reg93;
	        8'h5E   : reg_data_out <= slv_reg94;
	        8'h5F   : reg_data_out <= slv_reg95;
	        8'h60   : reg_data_out <= slv_reg96;
	        8'h61   : reg_data_out <= slv_reg97;
	        8'h62   : reg_data_out <= slv_reg98;
	        8'h63   : reg_data_out <= slv_reg99;
	        8'h64   : reg_data_out <= slv_reg100;
	        8'h65   : reg_data_out <= slv_reg101;
	        8'h66   : reg_data_out <= slv_reg102;
	        8'h67   : reg_data_out <= slv_reg103;
	        8'h68   : reg_data_out <= slv_reg104;
	        8'h69   : reg_data_out <= slv_reg105;
	        8'h6A   : reg_data_out <= slv_reg106;
	        8'h6B   : reg_data_out <= slv_reg107;
	        8'h6C   : reg_data_out <= slv_reg108;
	        8'h6D   : reg_data_out <= slv_reg109;
	        8'h6E   : reg_data_out <= slv_reg110;
	        8'h6F   : reg_data_out <= slv_reg111;
	        8'h70   : reg_data_out <= slv_reg112;
	        8'h71   : reg_data_out <= slv_reg113;
	        8'h72   : reg_data_out <= slv_reg114;
	        8'h73   : reg_data_out <= slv_reg115;
	        8'h74   : reg_data_out <= slv_reg116;
	        8'h75   : reg_data_out <= slv_reg117;
	        8'h76   : reg_data_out <= slv_reg118;
	        8'h77   : reg_data_out <= slv_reg119;
	        8'h78   : reg_data_out <= slv_reg120;
	        8'h79   : reg_data_out <= slv_reg121;
	        8'h7A   : reg_data_out <= slv_reg122;
	        8'h7B   : reg_data_out <= slv_reg123;
	        8'h7C   : reg_data_out <= slv_reg124;
	        8'h7D   : reg_data_out <= slv_reg125;
	        8'h7E   : reg_data_out <= slv_reg126;
	        8'h7F   : reg_data_out <= slv_reg127;
	        8'h80   : reg_data_out <= slv_reg128;
	        8'h81   : reg_data_out <= slv_reg129;
	        8'h82   : reg_data_out <= slv_reg130;
	        8'h83   : reg_data_out <= slv_reg131;
	        8'h84   : reg_data_out <= slv_reg132;
	        8'h85   : reg_data_out <= slv_reg133;
	        8'h86   : reg_data_out <= slv_reg134;
	        8'h87   : reg_data_out <= slv_reg135;
	        8'h88   : reg_data_out <= slv_reg136;
	        8'h89   : reg_data_out <= slv_reg137;
	        8'h8A   : reg_data_out <= slv_reg138;
	        8'h8B   : reg_data_out <= slv_reg139;
	        8'h8C   : reg_data_out <= slv_reg140;
	        8'h8D   : reg_data_out <= slv_reg141;
	        8'h8E   : reg_data_out <= slv_reg142;
	        8'h8F   : reg_data_out <= slv_reg143;
	        8'h90   : reg_data_out <= slv_reg144;
	        8'h91   : reg_data_out <= slv_reg145;
	        8'h92   : reg_data_out <= slv_reg146;
	        8'h93   : reg_data_out <= slv_reg147;
	        8'h94   : reg_data_out <= slv_reg148;
	        8'h95   : reg_data_out <= slv_reg149;
	        8'h96   : reg_data_out <= slv_reg150;
	        8'h97   : reg_data_out <= slv_reg151;
	        8'h98   : reg_data_out <= slv_reg152;
	        8'h99   : reg_data_out <= slv_reg153;
	        8'h9A   : reg_data_out <= slv_reg154;
	        8'h9B   : reg_data_out <= slv_reg155;
	        8'h9C   : reg_data_out <= slv_reg156;
	        8'h9D   : reg_data_out <= slv_reg157;
	        8'h9E   : reg_data_out <= slv_reg158;
	        8'h9F   : reg_data_out <= slv_reg159;
	        8'hA0   : reg_data_out <= slv_reg160;
	        8'hA1   : reg_data_out <= slv_reg161;
	        8'hA2   : reg_data_out <= slv_reg162;
	        8'hA3   : reg_data_out <= slv_reg163;
	        8'hA4   : reg_data_out <= slv_reg164;
	        8'hA5   : reg_data_out <= slv_reg165;
	        8'hA6   : reg_data_out <= slv_reg166;
	        8'hA7   : reg_data_out <= slv_reg167;
	        8'hA8   : reg_data_out <= slv_reg168;
	        8'hA9   : reg_data_out <= slv_reg169;
	        8'hAA   : reg_data_out <= slv_reg170;
	        8'hAB   : reg_data_out <= slv_reg171;
	        8'hAC   : reg_data_out <= slv_reg172;
	        8'hAD   : reg_data_out <= slv_reg173;
	        8'hAE   : reg_data_out <= slv_reg174;
	        8'hAF   : reg_data_out <= slv_reg175;
	        8'hB0   : reg_data_out <= slv_reg176;
	        8'hB1   : reg_data_out <= slv_reg177;
	        8'hB2   : reg_data_out <= slv_reg178;
	        8'hB3   : reg_data_out <= slv_reg179;
	        8'hB4   : reg_data_out <= slv_reg180;
	        8'hB5   : reg_data_out <= slv_reg181;
	        8'hB6   : reg_data_out <= slv_reg182;
	        8'hB7   : reg_data_out <= slv_reg183;
	        8'hB8   : reg_data_out <= slv_reg184;
	        8'hB9   : reg_data_out <= slv_reg185;
	        8'hBA   : reg_data_out <= slv_reg186;
	        8'hBB   : reg_data_out <= slv_reg187;
	        8'hBC   : reg_data_out <= slv_reg188;
	        8'hBD   : reg_data_out <= slv_reg189;
	        8'hBE   : reg_data_out <= slv_reg190;
	        8'hBF   : reg_data_out <= slv_reg191;
	        8'hC0   : reg_data_out <= slv_reg192;
	        8'hC1   : reg_data_out <= slv_reg193;
	        8'hC2   : reg_data_out <= slv_reg194;
	        8'hC3   : reg_data_out <= slv_reg195;
	        8'hC4   : reg_data_out <= slv_reg196;
	        8'hC5   : reg_data_out <= slv_reg197;
	        8'hC6   : reg_data_out <= slv_reg198;
	        8'hC7   : reg_data_out <= slv_reg199;
	        8'hC8   : reg_data_out <= slv_reg200;
	        8'hC9   : reg_data_out <= slv_reg201;
	        8'hCA   : reg_data_out <= slv_reg202;
	        8'hCB   : reg_data_out <= slv_reg203;
	        8'hCC   : reg_data_out <= slv_reg204;
	        8'hCD   : reg_data_out <= slv_reg205;
	        8'hCE   : reg_data_out <= slv_reg206;
	        8'hCF   : reg_data_out <= slv_reg207;
	        8'hD0   : reg_data_out <= slv_reg208;
	        8'hD1   : reg_data_out <= slv_reg209;
	        8'hD2   : reg_data_out <= slv_reg210;
	        8'hD3   : reg_data_out <= slv_reg211;
	        8'hD4   : reg_data_out <= slv_reg212;
	        8'hD5   : reg_data_out <= slv_reg213;
	        8'hD6   : reg_data_out <= slv_reg214;
	        8'hD7   : reg_data_out <= slv_reg215;
	        8'hD8   : reg_data_out <= slv_reg216;
	        8'hD9   : reg_data_out <= slv_reg217;
	        8'hDA   : reg_data_out <= slv_reg218;
	        8'hDB   : reg_data_out <= slv_reg219;
	        8'hDC   : reg_data_out <= slv_reg220;
	        8'hDD   : reg_data_out <= slv_reg221;
	        8'hDE   : reg_data_out <= slv_reg222;
	        8'hDF   : reg_data_out <= slv_reg223;
	        8'hE0   : reg_data_out <= slv_reg224;
	        8'hE1   : reg_data_out <= slv_reg225;
	        8'hE2   : reg_data_out <= slv_reg226;
	        8'hE3   : reg_data_out <= slv_reg227;
	        8'hE4   : reg_data_out <= slv_reg228;
	        8'hE5   : reg_data_out <= slv_reg229;
	        8'hE6   : reg_data_out <= slv_reg230;
	        8'hE7   : reg_data_out <= slv_reg231;
	        8'hE8   : reg_data_out <= slv_reg232;
	        8'hE9   : reg_data_out <= slv_reg233;
	        8'hEA   : reg_data_out <= slv_reg234;
	        8'hEB   : reg_data_out <= slv_reg235;
	        8'hEC   : reg_data_out <= slv_reg236;
	        8'hED   : reg_data_out <= slv_reg237;
	        8'hEE   : reg_data_out <= slv_reg238;
	        8'hEF   : reg_data_out <= slv_reg239;
	        8'hF0   : reg_data_out <= slv_reg240;
	        8'hF1   : reg_data_out <= slv_reg241;
	        8'hF2   : reg_data_out <= slv_reg242;
	        8'hF3   : reg_data_out <= slv_reg243;
	        8'hF4   : reg_data_out <= slv_reg244;
	        8'hF5   : reg_data_out <= slv_reg245;
	        8'hF6   : reg_data_out <= slv_reg246;
	        8'hF7   : reg_data_out <= slv_reg247;
	        8'hF8   : reg_data_out <= slv_reg248;
	        8'hF9   : reg_data_out <= slv_reg249;
	        8'hFA   : reg_data_out <= slv_reg250;
	        8'hFB   : reg_data_out <= slv_reg251;
	        8'hFC   : reg_data_out <= slv_reg252;
	        8'hFD   : reg_data_out <= slv_reg253;
	        8'hFE   : reg_data_out <= slv_reg254;
	        8'hFF   : reg_data_out <= slv_reg255;
            default : reg_data_out <= 0;
        endcase
	end

	always @(posedge S_AXI_ACLK) begin
        // Output register or memory read data
	    if(S_AXI_ARESETN == 1'b0) begin
	        axi_rdata  <= 0;
	    end
	    else begin
            // When there is a valid read address (S_AXI_ARVALID) with 
            // acceptance of read address by the slave (axi_arready), 
            // output the read dada 
            if(slv_reg_rden) begin
                axi_rdata <= reg_data_out;     // register read data
            end   
	    end
	end    

    // 2. RVALID & RRESP
    // axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both S_AXI_ARVALID and axi_arready are asserted.
    // The slave register's data are available on the axi_rdata bus at this instance.
    // The assertion of axi_rvalid marks the validity of read data on the bus and axi_rresp indicates the status of read transaction.
    // axi_rvalid is deasserted on reset (active low).
    // axi_rresp and axi_rdata are cleared to zero on reset (active low).
	always @(posedge S_AXI_ACLK) begin
        if(S_AXI_ARESETN == 1'b0) begin
            axi_rvalid <= 0;
            axi_rresp  <= 0;
	    end 
	    else begin
	        if(axi_arready && S_AXI_ARVALID && ~axi_rvalid) begin
                // Valid read data is available at the read data bus
                axi_rvalid <= 1'b1;
                axi_rresp  <= 2'b0; // 'OKAY' response
	        end   
	        else if(axi_rvalid && S_AXI_RREADY) begin
                // Read data is accepted by the master
                axi_rvalid <= 1'b0;
	        end                
	    end
	end

    // AXI4-Lite Interface Ends
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// Add User Custom Logic Here

// ============================================================================ //
//                                                                              //
//                                  Wire & Reg                                  //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Variable used for Core                                          //
// ==================================================================== //
    // 1. Variable for Input Registration
    // # User Guide : Comment the Registers which are Write Registers
    reg [31:0]  reg_64bit_1th_hi;
    reg [31:0]  reg_64bit_1th_lo;
    reg [31:0]  reg_64bit_2th_hi;
    reg [31:0]  reg_64bit_2th_lo;
    reg [31:0]  reg_64bit_3th_hi;
    reg [31:0]  reg_64bit_3th_lo;
    reg [31:0]  reg_64bit_4th_hi;
    reg [31:0]  reg_64bit_4th_lo;
    reg [31:0]  reg_64bit_5th_hi;
    reg [31:0]  reg_64bit_5th_lo;
    reg [31:0]  reg_64bit_6th_hi;
    reg [31:0]  reg_64bit_6th_lo;
    reg [31:0]  reg_64bit_7th_hi;
    reg [31:0]  reg_64bit_7th_lo;
    reg [31:0]  reg_64bit_8th_hi;
    reg [31:0]  reg_64bit_8th_lo;
    reg [31:0]  reg_64bit_9th_hi;
    reg [31:0]  reg_64bit_9th_lo;
    reg [31:0]  reg_64bit_10th_hi;
    reg [31:0]  reg_64bit_10th_lo;
    reg [31:0]  reg_64bit_11th_hi;
    reg [31:0]  reg_64bit_11th_lo;
    reg [31:0]  reg_64bit_12th_hi;
    reg [31:0]  reg_64bit_12th_lo;
    reg [31:0]  reg_64bit_13th_hi;
    reg [31:0]  reg_64bit_13th_lo;
    reg [31:0]  reg_64bit_14th_hi;
    reg [31:0]  reg_64bit_14th_lo;
    reg [31:0]  reg_64bit_15th_hi;
    reg [31:0]  reg_64bit_15th_lo;
    reg [31:0]  reg_64bit_16th_hi;
    reg [31:0]  reg_64bit_16th_lo;
    reg [31:0]  reg_64bit_17th_hi;
    reg [31:0]  reg_64bit_17th_lo;
    reg [31:0]  reg_64bit_18th_hi;
    reg [31:0]  reg_64bit_18th_lo;
    reg [31:0]  reg_64bit_19th_hi;
    reg [31:0]  reg_64bit_19th_lo;
    reg [31:0]  reg_64bit_20th_hi;
    reg [31:0]  reg_64bit_20th_lo;
    reg [31:0]  reg_64bit_21th_hi;
    reg [31:0]  reg_64bit_21th_lo;
    reg [31:0]  reg_64bit_22th_hi;
    reg [31:0]  reg_64bit_22th_lo;
    reg [31:0]  reg_64bit_23th_hi;
    reg [31:0]  reg_64bit_23th_lo;
    reg [31:0]  reg_64bit_24th_hi;
    reg [31:0]  reg_64bit_24th_lo;
    reg [31:0]  reg_64bit_25th_hi;
    reg [31:0]  reg_64bit_25th_lo;
    reg [31:0]  reg_64bit_26th_hi;
    reg [31:0]  reg_64bit_26th_lo;
    reg [31:0]  reg_64bit_27th_hi;
    reg [31:0]  reg_64bit_27th_lo;
    reg [31:0]  reg_64bit_28th_hi;
    reg [31:0]  reg_64bit_28th_lo;
    reg [31:0]  reg_64bit_29th_hi;
    reg [31:0]  reg_64bit_29th_lo;
    reg [31:0]  reg_64bit_30th_hi;
    reg [31:0]  reg_64bit_30th_lo;
    reg [31:0]  reg_64bit_31th_hi;
    reg [31:0]  reg_64bit_31th_lo;
    reg [31:0]  reg_64bit_32th_hi;
    reg [31:0]  reg_64bit_32th_lo;
    reg [31:0]  reg_64bit_33th_hi;
    reg [31:0]  reg_64bit_33th_lo;
    reg [31:0]  reg_64bit_34th_hi;
    reg [31:0]  reg_64bit_34th_lo;
    reg [31:0]  reg_64bit_35th_hi;
    reg [31:0]  reg_64bit_35th_lo;
    reg [31:0]  reg_64bit_36th_hi;
    reg [31:0]  reg_64bit_36th_lo;
    reg [31:0]  reg_64bit_37th_hi;
    reg [31:0]  reg_64bit_37th_lo;
    reg [31:0]  reg_64bit_38th_hi;
    reg [31:0]  reg_64bit_38th_lo;
    reg [31:0]  reg_64bit_39th_hi;
    reg [31:0]  reg_64bit_39th_lo;
    reg [31:0]  reg_64bit_40th_hi;
    reg [31:0]  reg_64bit_40th_lo;
    reg [31:0]  reg_64bit_41th_hi;
    reg [31:0]  reg_64bit_41th_lo;
    reg [31:0]  reg_64bit_42th_hi;
    reg [31:0]  reg_64bit_42th_lo;
    reg [31:0]  reg_64bit_43th_hi;
    reg [31:0]  reg_64bit_43th_lo;
    reg [31:0]  reg_64bit_44th_hi;
    reg [31:0]  reg_64bit_44th_lo;
    reg [31:0]  reg_64bit_45th_hi;
    reg [31:0]  reg_64bit_45th_lo;
    reg [31:0]  reg_64bit_46th_hi;
    reg [31:0]  reg_64bit_46th_lo;
    reg [31:0]  reg_64bit_47th_hi;
    reg [31:0]  reg_64bit_47th_lo;
    reg [31:0]  reg_64bit_48th_hi;
    reg [31:0]  reg_64bit_48th_lo;
    reg [31:0]  reg_64bit_49th_hi;
    reg [31:0]  reg_64bit_49th_lo;
    reg [31:0]  reg_64bit_50th_hi;
    reg [31:0]  reg_64bit_50th_lo;
    reg [31:0]  reg_64bit_51th_hi;
    reg [31:0]  reg_64bit_51th_lo;
    reg [31:0]  reg_64bit_52th_hi;
    reg [31:0]  reg_64bit_52th_lo;
    reg [31:0]  reg_64bit_53th_hi;
    reg [31:0]  reg_64bit_53th_lo;
    reg [31:0]  reg_64bit_54th_hi;
    reg [31:0]  reg_64bit_54th_lo;
    reg [31:0]  reg_64bit_55th_hi;
    reg [31:0]  reg_64bit_55th_lo;
    reg [31:0]  reg_64bit_56th_hi;
    reg [31:0]  reg_64bit_56th_lo;
    reg [31:0]  reg_64bit_57th_hi;
    reg [31:0]  reg_64bit_57th_lo;
    reg [31:0]  reg_64bit_58th_hi;
    reg [31:0]  reg_64bit_58th_lo;
    reg [31:0]  reg_64bit_59th_hi;
    reg [31:0]  reg_64bit_59th_lo;
    reg [31:0]  reg_64bit_60th_hi;
    reg [31:0]  reg_64bit_60th_lo;
    reg [31:0]  reg_64bit_61th_hi;
    reg [31:0]  reg_64bit_61th_lo;
    reg [31:0]  reg_64bit_62th_hi;
    reg [31:0]  reg_64bit_62th_lo;
    reg [31:0]  reg_64bit_63th_hi;
    reg [31:0]  reg_64bit_63th_lo;
    reg [31:0]  reg_64bit_64th_hi;
    reg [31:0]  reg_64bit_64th_lo;
    reg [31:0]  reg_64bit_65th_hi;
    reg [31:0]  reg_64bit_65th_lo;
    reg [31:0]  reg_64bit_66th_hi;
    reg [31:0]  reg_64bit_66th_lo;
    reg [31:0]  reg_64bit_67th_hi;
    reg [31:0]  reg_64bit_67th_lo;
    reg [31:0]  reg_64bit_68th_hi;
    reg [31:0]  reg_64bit_68th_lo;
    reg [31:0]  reg_64bit_69th_hi;
    reg [31:0]  reg_64bit_69th_lo;
    reg [31:0]  reg_64bit_70th_hi;
    reg [31:0]  reg_64bit_70th_lo;
    reg [31:0]  reg_64bit_71th_hi;
    reg [31:0]  reg_64bit_71th_lo;
    reg [31:0]  reg_64bit_72th_hi;
    reg [31:0]  reg_64bit_72th_lo;
    reg [31:0]  reg_64bit_73th_hi;
    reg [31:0]  reg_64bit_73th_lo;
    reg [31:0]  reg_64bit_74th_hi;
    reg [31:0]  reg_64bit_74th_lo;
    reg [31:0]  reg_64bit_75th_hi;
    reg [31:0]  reg_64bit_75th_lo;
    reg [31:0]  reg_64bit_76th_hi;
    reg [31:0]  reg_64bit_76th_lo;
    reg [31:0]  reg_64bit_77th_hi;
    reg [31:0]  reg_64bit_77th_lo;
    reg [31:0]  reg_64bit_78th_hi;
    reg [31:0]  reg_64bit_78th_lo;
    reg [31:0]  reg_64bit_79th_hi;
    reg [31:0]  reg_64bit_79th_lo;
    reg [31:0]  reg_64bit_80th_hi;
    reg [31:0]  reg_64bit_80th_lo;
    reg [31:0]  reg_64bit_81th_hi;
    reg [31:0]  reg_64bit_81th_lo;
    reg [31:0]  reg_64bit_82th_hi;
    reg [31:0]  reg_64bit_82th_lo;
    reg [31:0]  reg_64bit_83th_hi;
    reg [31:0]  reg_64bit_83th_lo;
    reg [31:0]  reg_64bit_84th_hi;
    reg [31:0]  reg_64bit_84th_lo;
    reg [31:0]  reg_64bit_85th_hi;
    reg [31:0]  reg_64bit_85th_lo;
    reg [31:0]  reg_64bit_86th_hi;
    reg [31:0]  reg_64bit_86th_lo;
    reg [31:0]  reg_64bit_87th_hi;
    reg [31:0]  reg_64bit_87th_lo;
    reg [31:0]  reg_64bit_88th_hi;
    reg [31:0]  reg_64bit_88th_lo;
    reg [31:0]  reg_64bit_89th_hi;
    reg [31:0]  reg_64bit_89th_lo;
    reg [31:0]  reg_64bit_90th_hi;
    reg [31:0]  reg_64bit_90th_lo;
    reg [31:0]  reg_64bit_91th_hi;
    reg [31:0]  reg_64bit_91th_lo;
    reg [31:0]  reg_64bit_92th_hi;
    reg [31:0]  reg_64bit_92th_lo;
    reg [31:0]  reg_64bit_93th_hi;
    reg [31:0]  reg_64bit_93th_lo;
    reg [31:0]  reg_64bit_94th_hi;
    reg [31:0]  reg_64bit_94th_lo;
    reg [31:0]  reg_64bit_95th_hi;
    reg [31:0]  reg_64bit_95th_lo;
    reg [31:0]  reg_64bit_96th_hi;
    reg [31:0]  reg_64bit_96th_lo;
    reg [31:0]  reg_64bit_97th_hi;
    reg [31:0]  reg_64bit_97th_lo;
    reg [31:0]  reg_64bit_98th_hi;
    reg [31:0]  reg_64bit_98th_lo;
    reg [31:0]  reg_64bit_99th_hi;
    reg [31:0]  reg_64bit_99th_lo;
    reg [31:0]  reg_64bit_100th_hi;
    reg [31:0]  reg_64bit_100th_lo;
    reg [31:0]  reg_64bit_101th_hi;
    reg [31:0]  reg_64bit_101th_lo;
    reg [31:0]  reg_64bit_102th_hi;
    reg [31:0]  reg_64bit_102th_lo;
    reg [31:0]  reg_64bit_103th_hi;
    reg [31:0]  reg_64bit_103th_lo;
    reg [31:0]  reg_64bit_104th_hi;
    reg [31:0]  reg_64bit_104th_lo;
    reg [31:0]  reg_64bit_105th_hi;
    reg [31:0]  reg_64bit_105th_lo;
    reg [31:0]  reg_64bit_106th_hi;
    reg [31:0]  reg_64bit_106th_lo;
    reg [31:0]  reg_64bit_107th_hi;
    reg [31:0]  reg_64bit_107th_lo;
    reg [31:0]  reg_64bit_108th_hi;
    reg [31:0]  reg_64bit_108th_lo;
    reg [31:0]  reg_64bit_109th_hi;
    reg [31:0]  reg_64bit_109th_lo;
    reg [31:0]  reg_64bit_110th_hi;
    reg [31:0]  reg_64bit_110th_lo;
    reg [31:0]  reg_64bit_111th_hi;
    reg [31:0]  reg_64bit_111th_lo;
    reg [31:0]  reg_64bit_112th_hi;
    reg [31:0]  reg_64bit_112th_lo;
    reg [31:0]  reg_64bit_113th_hi;
    reg [31:0]  reg_64bit_113th_lo;
    reg [31:0]  reg_64bit_114th_hi;
    reg [31:0]  reg_64bit_114th_lo;
    reg [31:0]  reg_64bit_115th_hi;
    reg [31:0]  reg_64bit_115th_lo;
    reg [31:0]  reg_64bit_116th_hi;
    reg [31:0]  reg_64bit_116th_lo;
    reg [31:0]  reg_64bit_117th_hi;
    reg [31:0]  reg_64bit_117th_lo;
    reg [31:0]  reg_64bit_118th_hi;
    reg [31:0]  reg_64bit_118th_lo;
    reg [31:0]  reg_64bit_119th_hi;
    reg [31:0]  reg_64bit_119th_lo;
    reg [31:0]  reg_64bit_120th_hi;
    reg [31:0]  reg_64bit_120th_lo;
    reg [31:0]  reg_64bit_121th_hi;
    reg [31:0]  reg_64bit_121th_lo;
    reg [31:0]  reg_64bit_122th_hi;
    reg [31:0]  reg_64bit_122th_lo;
    reg [31:0]  reg_64bit_123th_hi;
    reg [31:0]  reg_64bit_123th_lo;
    reg [31:0]  reg_64bit_124th_hi;
    reg [31:0]  reg_64bit_124th_lo;
    reg [31:0]  reg_64bit_125th_hi;
    reg [31:0]  reg_64bit_125th_lo;
    reg [31:0]  reg_64bit_126th_hi;
    reg [31:0]  reg_64bit_126th_lo;
    reg [31:0]  reg_64bit_127th_hi;
    reg [31:0]  reg_64bit_127th_lo;
    reg [31:0]  reg_64bit_128th_hi;
    reg [31:0]  reg_64bit_128th_lo;

    // 2. Variable for Intermediate Process
    reg         upper_flag;
    reg [63:0]  captured_data;


// ============================================================================ //
//                                                                              //
//                                Input Regist.                                 //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Registration of Input Signals                                   //
// ==================================================================== //
    // # User Guide : Comment the Registers which are Write or Un-Used Registers
    // 1. 1st 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_1th_hi <= 0;
        else                    reg_64bit_1th_hi <= i_reg_64bit_1th_hi;
    end

    // 2. 1st 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_1th_lo <= 0;
        else                    reg_64bit_1th_lo <= i_reg_64bit_1th_lo;
    end

    // 3. 2nd 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_2th_hi <= 0;
        else                    reg_64bit_2th_hi <= i_reg_64bit_2th_hi;
    end

    // 4. 2nd 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_2th_lo <= 0;
        else                    reg_64bit_2th_lo <= i_reg_64bit_2th_lo;
    end

    // 5. 3th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_3th_hi <= 0;
        else                    reg_64bit_3th_hi <= i_reg_64bit_3th_hi;
    end

    // 6. 3th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_3th_lo <= 0;
        else                    reg_64bit_3th_lo <= i_reg_64bit_3th_lo;
    end

    // 7. 4th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_4th_hi <= 0;
        else                    reg_64bit_4th_hi <= i_reg_64bit_4th_hi;
    end

    // 8. 4th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_4th_lo <= 0;
        else                    reg_64bit_4th_lo <= i_reg_64bit_4th_lo;
    end

    // 9. 5th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_5th_hi <= 0;
        else                    reg_64bit_5th_hi <= i_reg_64bit_5th_hi;
    end

    // 10. 5th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_5th_lo <= 0;
        else                    reg_64bit_5th_lo <= i_reg_64bit_5th_lo;
    end

    // 11. 6th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_6th_hi <= 0;
        else                    reg_64bit_6th_hi <= i_reg_64bit_6th_hi;
    end

    // 12. 6th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_6th_lo <= 0;
        else                    reg_64bit_6th_lo <= i_reg_64bit_6th_lo;
    end

    // 13. 7th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_7th_hi <= 0;
        else                    reg_64bit_7th_hi <= i_reg_64bit_7th_hi;
    end

    // 14. 7th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_7th_lo <= 0;
        else                    reg_64bit_7th_lo <= i_reg_64bit_7th_lo;
    end

    // 15. 8th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_8th_hi <= 0;
        else                    reg_64bit_8th_hi <= i_reg_64bit_8th_hi;
    end

    // 16. 8th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_8th_lo <= 0;
        else                    reg_64bit_8th_lo <= i_reg_64bit_8th_lo;
    end

    // 17. 9th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_9th_hi <= 0;
        else                    reg_64bit_9th_hi <= i_reg_64bit_9th_hi;
    end

    // 18. 9th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_9th_lo <= 0;
        else                    reg_64bit_9th_lo <= i_reg_64bit_9th_lo;
    end

    // 19. 10th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_10th_hi <= 0;
        else                    reg_64bit_10th_hi <= i_reg_64bit_10th_hi;
    end

    // 20. 10th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_10th_lo <= 0;
        else                    reg_64bit_10th_lo <= i_reg_64bit_10th_lo;
    end

    // 21. 11th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_11th_hi <= 0;
        else                    reg_64bit_11th_hi <= i_reg_64bit_11th_hi;
    end

    // 22. 11th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_11th_lo <= 0;
        else                    reg_64bit_11th_lo <= i_reg_64bit_11th_lo;
    end

    // 23. 12th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_12th_hi <= 0;
        else                    reg_64bit_12th_hi <= i_reg_64bit_12th_hi;
    end

    // 24. 12th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_12th_lo <= 0;
        else                    reg_64bit_12th_lo <= i_reg_64bit_12th_lo;
    end

    // 25. 13th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_13th_hi <= 0;
        else                    reg_64bit_13th_hi <= i_reg_64bit_13th_hi;
    end

    // 26. 13th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_13th_lo <= 0;
        else                    reg_64bit_13th_lo <= i_reg_64bit_13th_lo;
    end

    // 27. 14th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_14th_hi <= 0;
        else                    reg_64bit_14th_hi <= i_reg_64bit_14th_hi;
    end

    // 28. 14th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_14th_lo <= 0;
        else                    reg_64bit_14th_lo <= i_reg_64bit_14th_lo;
    end

    // 29. 15th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_15th_hi <= 0;
        else                    reg_64bit_15th_hi <= i_reg_64bit_15th_hi;
    end

    // 30. 15th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_15th_lo <= 0;
        else                    reg_64bit_15th_lo <= i_reg_64bit_15th_lo;
    end

    // 31. 16th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_16th_hi <= 0;
        else                    reg_64bit_16th_hi <= i_reg_64bit_16th_hi;
    end

    // 32. 16th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_16th_lo <= 0;
        else                    reg_64bit_16th_lo <= i_reg_64bit_16th_lo;
    end

    // 33. 17th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_17th_hi <= 0;
        else                    reg_64bit_17th_hi <= i_reg_64bit_17th_hi;
    end

    // 34. 17th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_17th_lo <= 0;
        else                    reg_64bit_17th_lo <= i_reg_64bit_17th_lo;
    end

    // 35. 18th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_18th_hi <= 0;
        else                    reg_64bit_18th_hi <= i_reg_64bit_18th_hi;
    end

    // 36. 18th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_18th_lo <= 0;
        else                    reg_64bit_18th_lo <= i_reg_64bit_18th_lo;
    end

    // 37. 19th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_19th_hi <= 0;
        else                    reg_64bit_19th_hi <= i_reg_64bit_19th_hi;
    end

    // 38. 19th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_19th_lo <= 0;
        else                    reg_64bit_19th_lo <= i_reg_64bit_19th_lo;
    end

    // 39. 20th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_20th_hi <= 0;
        else                    reg_64bit_20th_hi <= i_reg_64bit_20th_hi;
    end

    // 40. 20th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_20th_lo <= 0;
        else                    reg_64bit_20th_lo <= i_reg_64bit_20th_lo;
    end

    // 41. 21th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_21th_hi <= 0;
        else                    reg_64bit_21th_hi <= i_reg_64bit_21th_hi;
    end

    // 42. 21th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_21th_lo <= 0;
        else                    reg_64bit_21th_lo <= i_reg_64bit_21th_lo;
    end

    // 43. 22th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_22th_hi <= 0;
        else                    reg_64bit_22th_hi <= i_reg_64bit_22th_hi;
    end

    // 44. 22th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_22th_lo <= 0;
        else                    reg_64bit_22th_lo <= i_reg_64bit_22th_lo;
    end

    // 45. 23th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_23th_hi <= 0;
        else                    reg_64bit_23th_hi <= i_reg_64bit_23th_hi;
    end

    // 46. 23th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_23th_lo <= 0;
        else                    reg_64bit_23th_lo <= i_reg_64bit_23th_lo;
    end

    // 47. 24th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_24th_hi <= 0;
        else                    reg_64bit_24th_hi <= i_reg_64bit_24th_hi;
    end

    // 48. 24th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_24th_lo <= 0;
        else                    reg_64bit_24th_lo <= i_reg_64bit_24th_lo;
    end

    // 49. 25th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_25th_hi <= 0;
        else                    reg_64bit_25th_hi <= i_reg_64bit_25th_hi;
    end

    // 50. 25th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_25th_lo <= 0;
        else                    reg_64bit_25th_lo <= i_reg_64bit_25th_lo;
    end

    // 51. 26th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_26th_hi <= 0;
        else                    reg_64bit_26th_hi <= i_reg_64bit_26th_hi;
    end

    // 52. 26th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_26th_lo <= 0;
        else                    reg_64bit_26th_lo <= i_reg_64bit_26th_lo;
    end

    // 53. 27th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_27th_hi <= 0;
        else                    reg_64bit_27th_hi <= i_reg_64bit_27th_hi;
    end

    // 54. 27th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_27th_lo <= 0;
        else                    reg_64bit_27th_lo <= i_reg_64bit_27th_lo;
    end

    // 55. 28th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_28th_hi <= 0;
        else                    reg_64bit_28th_hi <= i_reg_64bit_28th_hi;
    end

    // 56. 28th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_28th_lo <= 0;
        else                    reg_64bit_28th_lo <= i_reg_64bit_28th_lo;
    end

    // 57. 29th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_29th_hi <= 0;
        else                    reg_64bit_29th_hi <= i_reg_64bit_29th_hi;
    end

    // 58. 29th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_29th_lo <= 0;
        else                    reg_64bit_29th_lo <= i_reg_64bit_29th_lo;
    end

    // 59. 30th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_30th_hi <= 0;
        else                    reg_64bit_30th_hi <= i_reg_64bit_30th_hi;
    end

    // 60. 30th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_30th_lo <= 0;
        else                    reg_64bit_30th_lo <= i_reg_64bit_30th_lo;
    end

    // 61. 31th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_31th_hi <= 0;
        else                    reg_64bit_31th_hi <= i_reg_64bit_31th_hi;
    end

    // 62. 31th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_31th_lo <= 0;
        else                    reg_64bit_31th_lo <= i_reg_64bit_31th_lo;
    end

    // 63. 32th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_32th_hi <= 0;
        else                    reg_64bit_32th_hi <= i_reg_64bit_32th_hi;
    end

    // 64. 32th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_32th_lo <= 0;
        else                    reg_64bit_32th_lo <= i_reg_64bit_32th_lo;
    end

    // 65. 33th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_33th_hi <= 0;
        else                    reg_64bit_33th_hi <= i_reg_64bit_33th_hi;
    end

    // 66. 33th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_33th_lo <= 0;
        else                    reg_64bit_33th_lo <= i_reg_64bit_33th_lo;
    end

    // 67. 34th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_34th_hi <= 0;
        else                    reg_64bit_34th_hi <= i_reg_64bit_34th_hi;
    end

    // 68. 34th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_34th_lo <= 0;
        else                    reg_64bit_34th_lo <= i_reg_64bit_34th_lo;
    end

    // 69. 35th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_35th_hi <= 0;
        else                    reg_64bit_35th_hi <= i_reg_64bit_35th_hi;
    end

    // 70. 35th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_35th_lo <= 0;
        else                    reg_64bit_35th_lo <= i_reg_64bit_35th_lo;
    end

    // 71. 36th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_36th_hi <= 0;
        else                    reg_64bit_36th_hi <= i_reg_64bit_36th_hi;
    end

    // 72. 36th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_36th_lo <= 0;
        else                    reg_64bit_36th_lo <= i_reg_64bit_36th_lo;
    end

    // 73. 37th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_37th_hi <= 0;
        else                    reg_64bit_37th_hi <= i_reg_64bit_37th_hi;
    end

    // 74. 37th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_37th_lo <= 0;
        else                    reg_64bit_37th_lo <= i_reg_64bit_37th_lo;
    end

    // 75. 38th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_38th_hi <= 0;
        else                    reg_64bit_38th_hi <= i_reg_64bit_38th_hi;
    end

    // 76. 38th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_38th_lo <= 0;
        else                    reg_64bit_38th_lo <= i_reg_64bit_38th_lo;
    end

    // 77. 39th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_39th_hi <= 0;
        else                    reg_64bit_39th_hi <= i_reg_64bit_39th_hi;
    end

    // 78. 39th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_39th_lo <= 0;
        else                    reg_64bit_39th_lo <= i_reg_64bit_39th_lo;
    end

    // 79. 40th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_40th_hi <= 0;
        else                    reg_64bit_40th_hi <= i_reg_64bit_40th_hi;
    end

    // 80. 40th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_40th_lo <= 0;
        else                    reg_64bit_40th_lo <= i_reg_64bit_40th_lo;
    end

    // 81. 41th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_41th_hi <= 0;
        else                    reg_64bit_41th_hi <= i_reg_64bit_41th_hi;
    end

    // 82. 41th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_41th_lo <= 0;
        else                    reg_64bit_41th_lo <= i_reg_64bit_41th_lo;
    end

    // 83. 42th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_42th_hi <= 0;
        else                    reg_64bit_42th_hi <= i_reg_64bit_42th_hi;
    end

    // 84. 42th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_42th_lo <= 0;
        else                    reg_64bit_42th_lo <= i_reg_64bit_42th_lo;
    end

    // 85. 43th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_43th_hi <= 0;
        else                    reg_64bit_43th_hi <= i_reg_64bit_43th_hi;
    end

    // 86. 43th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_43th_lo <= 0;
        else                    reg_64bit_43th_lo <= i_reg_64bit_43th_lo;
    end

    // 87. 44th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_44th_hi <= 0;
        else                    reg_64bit_44th_hi <= i_reg_64bit_44th_hi;
    end

    // 88. 44th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_44th_lo <= 0;
        else                    reg_64bit_44th_lo <= i_reg_64bit_44th_lo;
    end

    // 89. 45th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_45th_hi <= 0;
        else                    reg_64bit_45th_hi <= i_reg_64bit_45th_hi;
    end

    // 90. 45th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_45th_lo <= 0;
        else                    reg_64bit_45th_lo <= i_reg_64bit_45th_lo;
    end

    // 91. 46th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_46th_hi <= 0;
        else                    reg_64bit_46th_hi <= i_reg_64bit_46th_hi;
    end

    // 92. 46th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_46th_lo <= 0;
        else                    reg_64bit_46th_lo <= i_reg_64bit_46th_lo;
    end

    // 93. 47th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_47th_hi <= 0;
        else                    reg_64bit_47th_hi <= i_reg_64bit_47th_hi;
    end

    // 94. 47th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_47th_lo <= 0;
        else                    reg_64bit_47th_lo <= i_reg_64bit_47th_lo;
    end

    // 95. 48th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_48th_hi <= 0;
        else                    reg_64bit_48th_hi <= i_reg_64bit_48th_hi;
    end

    // 96. 48th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_48th_lo <= 0;
        else                    reg_64bit_48th_lo <= i_reg_64bit_48th_lo;
    end

    // 97. 49th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_49th_hi <= 0;
        else                    reg_64bit_49th_hi <= i_reg_64bit_49th_hi;
    end

    // 98. 49th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_49th_lo <= 0;
        else                    reg_64bit_49th_lo <= i_reg_64bit_49th_lo;
    end

    // 99. 50th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_50th_hi <= 0;
        else                    reg_64bit_50th_hi <= i_reg_64bit_50th_hi;
    end

    // 100. 50th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_50th_lo <= 0;
        else                    reg_64bit_50th_lo <= i_reg_64bit_50th_lo;
    end

    // 101. 51th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_51th_hi <= 0;
        else                    reg_64bit_51th_hi <= i_reg_64bit_51th_hi;
    end

    // 102. 51th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_51th_lo <= 0;
        else                    reg_64bit_51th_lo <= i_reg_64bit_51th_lo;
    end

    // 103. 52th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_52th_hi <= 0;
        else                    reg_64bit_52th_hi <= i_reg_64bit_52th_hi;
    end

    // 104. 52th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_52th_lo <= 0;
        else                    reg_64bit_52th_lo <= i_reg_64bit_52th_lo;
    end

    // 105. 53th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_53th_hi <= 0;
        else                    reg_64bit_53th_hi <= i_reg_64bit_53th_hi;
    end

    // 106. 53th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_53th_lo <= 0;
        else                    reg_64bit_53th_lo <= i_reg_64bit_53th_lo;
    end

    // 107. 54th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_54th_hi <= 0;
        else                    reg_64bit_54th_hi <= i_reg_64bit_54th_hi;
    end

    // 108. 54th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_54th_lo <= 0;
        else                    reg_64bit_54th_lo <= i_reg_64bit_54th_lo;
    end

    // 109. 55th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_55th_hi <= 0;
        else                    reg_64bit_55th_hi <= i_reg_64bit_55th_hi;
    end

    // 110. 55th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_55th_lo <= 0;
        else                    reg_64bit_55th_lo <= i_reg_64bit_55th_lo;
    end

    // 111. 56th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_56th_hi <= 0;
        else                    reg_64bit_56th_hi <= i_reg_64bit_56th_hi;
    end

    // 112. 56th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_56th_lo <= 0;
        else                    reg_64bit_56th_lo <= i_reg_64bit_56th_lo;
    end

    // 113. 57th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_57th_hi <= 0;
        else                    reg_64bit_57th_hi <= i_reg_64bit_57th_hi;
    end

    // 114. 57th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_57th_lo <= 0;
        else                    reg_64bit_57th_lo <= i_reg_64bit_57th_lo;
    end

    // 115. 58th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_58th_hi <= 0;
        else                    reg_64bit_58th_hi <= i_reg_64bit_58th_hi;
    end

    // 116. 58th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_58th_lo <= 0;
        else                    reg_64bit_58th_lo <= i_reg_64bit_58th_lo;
    end

    // 117. 59th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_59th_hi <= 0;
        else                    reg_64bit_59th_hi <= i_reg_64bit_59th_hi;
    end

    // 118. 59th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_59th_lo <= 0;
        else                    reg_64bit_59th_lo <= i_reg_64bit_59th_lo;
    end

    // 119. 60th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_60th_hi <= 0;
        else                    reg_64bit_60th_hi <= i_reg_64bit_60th_hi;
    end

    // 120. 60th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_60th_lo <= 0;
        else                    reg_64bit_60th_lo <= i_reg_64bit_60th_lo;
    end

    // 121. 61th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_61th_hi <= 0;
        else                    reg_64bit_61th_hi <= i_reg_64bit_61th_hi;
    end

    // 122. 61th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_61th_lo <= 0;
        else                    reg_64bit_61th_lo <= i_reg_64bit_61th_lo;
    end

    // 123. 62th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_62th_hi <= 0;
        else                    reg_64bit_62th_hi <= i_reg_64bit_62th_hi;
    end

    // 124. 62th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_62th_lo <= 0;
        else                    reg_64bit_62th_lo <= i_reg_64bit_62th_lo;
    end

    // 125. 63th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_63th_hi <= 0;
        else                    reg_64bit_63th_hi <= i_reg_64bit_63th_hi;
    end

    // 126. 63th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_63th_lo <= 0;
        else                    reg_64bit_63th_lo <= i_reg_64bit_63th_lo;
    end

    // 127. 64th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_64th_hi <= 0;
        else                    reg_64bit_64th_hi <= i_reg_64bit_64th_hi;
    end

    // 128. 64th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_64th_lo <= 0;
        else                    reg_64bit_64th_lo <= i_reg_64bit_64th_lo;
    end

    // 129. 65th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_65th_hi <= 0;
        else                    reg_64bit_65th_hi <= i_reg_64bit_65th_hi;
    end

    // 130. 65th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_65th_lo <= 0;
        else                    reg_64bit_65th_lo <= i_reg_64bit_65th_lo;
    end

    // 131. 66th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_66th_hi <= 0;
        else                    reg_64bit_66th_hi <= i_reg_64bit_66th_hi;
    end

    // 132. 66th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_66th_lo <= 0;
        else                    reg_64bit_66th_lo <= i_reg_64bit_66th_lo;
    end

    // 133. 67th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_67th_hi <= 0;
        else                    reg_64bit_67th_hi <= i_reg_64bit_67th_hi;
    end

    // 134. 67th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_67th_lo <= 0;
        else                    reg_64bit_67th_lo <= i_reg_64bit_67th_lo;
    end

    // 135. 68th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_68th_hi <= 0;
        else                    reg_64bit_68th_hi <= i_reg_64bit_68th_hi;
    end

    // 136. 68th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_68th_lo <= 0;
        else                    reg_64bit_68th_lo <= i_reg_64bit_68th_lo;
    end

    // 137. 69th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_69th_hi <= 0;
        else                    reg_64bit_69th_hi <= i_reg_64bit_69th_hi;
    end

    // 138. 69th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_69th_lo <= 0;
        else                    reg_64bit_69th_lo <= i_reg_64bit_69th_lo;
    end

    // 139. 70th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_70th_hi <= 0;
        else                    reg_64bit_70th_hi <= i_reg_64bit_70th_hi;
    end

    // 140. 70th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_70th_lo <= 0;
        else                    reg_64bit_70th_lo <= i_reg_64bit_70th_lo;
    end

    // 141. 71th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_71th_hi <= 0;
        else                    reg_64bit_71th_hi <= i_reg_64bit_71th_hi;
    end

    // 142. 71th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_71th_lo <= 0;
        else                    reg_64bit_71th_lo <= i_reg_64bit_71th_lo;
    end

    // 143. 72th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_72th_hi <= 0;
        else                    reg_64bit_72th_hi <= i_reg_64bit_72th_hi;
    end

    // 144. 72th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_72th_lo <= 0;
        else                    reg_64bit_72th_lo <= i_reg_64bit_72th_lo;
    end

    // 145. 73th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_73th_hi <= 0;
        else                    reg_64bit_73th_hi <= i_reg_64bit_73th_hi;
    end

    // 146. 73th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_73th_lo <= 0;
        else                    reg_64bit_73th_lo <= i_reg_64bit_73th_lo;
    end

    // 147. 74th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_74th_hi <= 0;
        else                    reg_64bit_74th_hi <= i_reg_64bit_74th_hi;
    end

    // 148. 74th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_74th_lo <= 0;
        else                    reg_64bit_74th_lo <= i_reg_64bit_74th_lo;
    end
    
    // 149. 75th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_75th_hi <= 0;
        else                    reg_64bit_75th_hi <= i_reg_64bit_75th_hi;
    end

    // 150. 75th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_75th_lo <= 0;
        else                    reg_64bit_75th_lo <= i_reg_64bit_75th_lo;
    end

    // 151. 76th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_76th_hi <= 0;
        else                    reg_64bit_76th_hi <= i_reg_64bit_76th_hi;
    end

    // 152. 76th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_76th_lo <= 0;
        else                    reg_64bit_76th_lo <= i_reg_64bit_76th_lo;
    end

    // 153. 77th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_77th_hi <= 0;
        else                    reg_64bit_77th_hi <= i_reg_64bit_77th_hi;
    end

    // 154. 77th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_77th_lo <= 0;
        else                    reg_64bit_77th_lo <= i_reg_64bit_77th_lo;
    end

    // 155. 78th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_78th_hi <= 0;
        else                    reg_64bit_78th_hi <= i_reg_64bit_78th_hi;
    end

    // 156. 78th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_78th_lo <= 0;
        else                    reg_64bit_78th_lo <= i_reg_64bit_78th_lo;
    end

    // 157. 79th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_79th_hi <= 0;
        else                    reg_64bit_79th_hi <= i_reg_64bit_79th_hi;
    end

    // 158. 79th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_79th_lo <= 0;
        else                    reg_64bit_79th_lo <= i_reg_64bit_79th_lo;
    end

    // 159. 80th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_80th_hi <= 0;
        else                    reg_64bit_80th_hi <= i_reg_64bit_80th_hi;
    end

    // 160. 80th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_80th_lo <= 0;
        else                    reg_64bit_80th_lo <= i_reg_64bit_80th_lo;
    end

    // 161. 81th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_81th_hi <= 0;
        else                    reg_64bit_81th_hi <= i_reg_64bit_81th_hi;
    end

    // 162. 81th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_81th_lo <= 0;
        else                    reg_64bit_81th_lo <= i_reg_64bit_81th_lo;
    end

    // 163. 82th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_82th_hi <= 0;
        else                    reg_64bit_82th_hi <= i_reg_64bit_82th_hi;
    end

    // 164. 82th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_82th_lo <= 0;
        else                    reg_64bit_82th_lo <= i_reg_64bit_82th_lo;
    end

    // 165. 83th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_83th_hi <= 0;
        else                    reg_64bit_83th_hi <= i_reg_64bit_83th_hi;
    end

    // 166. 83th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_83th_lo <= 0;
        else                    reg_64bit_83th_lo <= i_reg_64bit_83th_lo;
    end

    // 167. 84th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_84th_hi <= 0;
        else                    reg_64bit_84th_hi <= i_reg_64bit_84th_hi;
    end

    // 168. 84th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_84th_lo <= 0;
        else                    reg_64bit_84th_lo <= i_reg_64bit_84th_lo;
    end

    // 169. 85th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_85th_hi <= 0;
        else                    reg_64bit_85th_hi <= i_reg_64bit_85th_hi;
    end

    // 170. 85th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_85th_lo <= 0;
        else                    reg_64bit_85th_lo <= i_reg_64bit_85th_lo;
    end

    // 171. 86th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_86th_hi <= 0;
        else                    reg_64bit_86th_hi <= i_reg_64bit_86th_hi;
    end

    // 172. 86th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_86th_lo <= 0;
        else                    reg_64bit_86th_lo <= i_reg_64bit_86th_lo;
    end

    // 173. 87th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_87th_hi <= 0;
        else                    reg_64bit_87th_hi <= i_reg_64bit_87th_hi;
    end

    // 174. 87th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_87th_lo <= 0;
        else                    reg_64bit_87th_lo <= i_reg_64bit_87th_lo;
    end

    // 175. 88th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_88th_hi <= 0;
        else                    reg_64bit_88th_hi <= i_reg_64bit_88th_hi;
    end

    // 176. 88th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_88th_lo <= 0;
        else                    reg_64bit_88th_lo <= i_reg_64bit_88th_lo;
    end

    // 177. 89th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_89th_hi <= 0;
        else                    reg_64bit_89th_hi <= i_reg_64bit_89th_hi;
    end

    // 178. 89th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_89th_lo <= 0;
        else                    reg_64bit_89th_lo <= i_reg_64bit_89th_lo;
    end

    // 179. 90th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_90th_hi <= 0;
        else                    reg_64bit_90th_hi <= i_reg_64bit_90th_hi;
    end

    // 180. 90th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_90th_lo <= 0;
        else                    reg_64bit_90th_lo <= i_reg_64bit_90th_lo;
    end

    // 181. 91th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_91th_hi <= 0;
        else                    reg_64bit_91th_hi <= i_reg_64bit_91th_hi;
    end

    // 182. 91th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_91th_lo <= 0;
        else                    reg_64bit_91th_lo <= i_reg_64bit_91th_lo;
    end

    // 183. 92th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_92th_hi <= 0;
        else                    reg_64bit_92th_hi <= i_reg_64bit_92th_hi;
    end

    // 184. 92th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_92th_lo <= 0;
        else                    reg_64bit_92th_lo <= i_reg_64bit_92th_lo;
    end

    // 185. 93th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_93th_hi <= 0;
        else                    reg_64bit_93th_hi <= i_reg_64bit_93th_hi;
    end

    // 186. 93th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_93th_lo <= 0;
        else                    reg_64bit_93th_lo <= i_reg_64bit_93th_lo;
    end

    // 187. 94th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_94th_hi <= 0;
        else                    reg_64bit_94th_hi <= i_reg_64bit_94th_hi;
    end

    // 188. 94th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_94th_lo <= 0;
        else                    reg_64bit_94th_lo <= i_reg_64bit_94th_lo;
    end

    // 189. 95th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_95th_hi <= 0;
        else                    reg_64bit_95th_hi <= i_reg_64bit_95th_hi;
    end

    // 190. 95th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_95th_lo <= 0;
        else                    reg_64bit_95th_lo <= i_reg_64bit_95th_lo;
    end

    // 191. 96th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_96th_hi <= 0;
        else                    reg_64bit_96th_hi <= i_reg_64bit_96th_hi;
    end

    // 192. 96th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_96th_lo <= 0;
        else                    reg_64bit_96th_lo <= i_reg_64bit_96th_lo;
    end

    // 193. 97th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_97th_hi <= 0;
        else                    reg_64bit_97th_hi <= i_reg_64bit_97th_hi;
    end

    // 194. 97th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_97th_lo <= 0;
        else                    reg_64bit_97th_lo <= i_reg_64bit_97th_lo;
    end

    // 195. 98th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_98th_hi <= 0;
        else                    reg_64bit_98th_hi <= i_reg_64bit_98th_hi;
    end

    // 196. 98th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_98th_lo <= 0;
        else                    reg_64bit_98th_lo <= i_reg_64bit_98th_lo;
    end

    // 197. 99th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_99th_hi <= 0;
        else                    reg_64bit_99th_hi <= i_reg_64bit_99th_hi;
    end

    // 198. 99th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_99th_lo <= 0;
        else                    reg_64bit_99th_lo <= i_reg_64bit_99th_lo;
    end

    // 199. 100th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_100th_hi <= 0;
        else                    reg_64bit_100th_hi <= i_reg_64bit_100th_hi;
    end

    // 200. 100th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_100th_lo <= 0;
        else                    reg_64bit_100th_lo <= i_reg_64bit_100th_lo;
    end

    // 201. 101th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_101th_hi <= 0;
        else                    reg_64bit_101th_hi <= i_reg_64bit_101th_hi;
    end

    // 202. 101th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_101th_lo <= 0;
        else                    reg_64bit_101th_lo <= i_reg_64bit_101th_lo;
    end

    // 203. 102th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_102th_hi <= 0;
        else                    reg_64bit_102th_hi <= i_reg_64bit_102th_hi;
    end

    // 204. 102th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_102th_lo <= 0;
        else                    reg_64bit_102th_lo <= i_reg_64bit_102th_lo;
    end

    // 205. 103th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_103th_hi <= 0;
        else                    reg_64bit_103th_hi <= i_reg_64bit_103th_hi;
    end

    // 206. 103th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_103th_lo <= 0;
        else                    reg_64bit_103th_lo <= i_reg_64bit_103th_lo;
    end

    // 207. 104th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_104th_hi <= 0;
        else                    reg_64bit_104th_hi <= i_reg_64bit_104th_hi;
    end

    // 208. 104th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_104th_lo <= 0;
        else                    reg_64bit_104th_lo <= i_reg_64bit_104th_lo;
    end

    // 209. 105th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_105th_hi <= 0;
        else                    reg_64bit_105th_hi <= i_reg_64bit_105th_hi;
    end

    // 210. 105th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_105th_lo <= 0;
        else                    reg_64bit_105th_lo <= i_reg_64bit_105th_lo;
    end

    // 211. 106th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_106th_hi <= 0;
        else                    reg_64bit_106th_hi <= i_reg_64bit_106th_hi;
    end

    // 212. 106th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_106th_lo <= 0;
        else                    reg_64bit_106th_lo <= i_reg_64bit_106th_lo;
    end

    // 213. 107th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_107th_hi <= 0;
        else                    reg_64bit_107th_hi <= i_reg_64bit_107th_hi;
    end

    // 214. 107th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_107th_lo <= 0;
        else                    reg_64bit_107th_lo <= i_reg_64bit_107th_lo;
    end

    // 215. 108th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_108th_hi <= 0;
        else                    reg_64bit_108th_hi <= i_reg_64bit_108th_hi;
    end

    // 216. 108th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_108th_lo <= 0;
        else                    reg_64bit_108th_lo <= i_reg_64bit_108th_lo;
    end

    // 217. 109th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_109th_hi <= 0;
        else                    reg_64bit_109th_hi <= i_reg_64bit_109th_hi;
    end

    // 218. 109th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_109th_lo <= 0;
        else                    reg_64bit_109th_lo <= i_reg_64bit_109th_lo;
    end

    // 219. 110th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_110th_hi <= 0;
        else                    reg_64bit_110th_hi <= i_reg_64bit_110th_hi;
    end

    // 220. 110th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_110th_lo <= 0;
        else                    reg_64bit_110th_lo <= i_reg_64bit_110th_lo;
    end

    // 221. 111th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_111th_hi <= 0;
        else                    reg_64bit_111th_hi <= i_reg_64bit_111th_hi;
    end

    // 222. 111th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_111th_lo <= 0;
        else                    reg_64bit_111th_lo <= i_reg_64bit_111th_lo;
    end

    // 223. 112th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_112th_hi <= 0;
        else                    reg_64bit_112th_hi <= i_reg_64bit_112th_hi;
    end

    // 224. 112th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_112th_lo <= 0;
        else                    reg_64bit_112th_lo <= i_reg_64bit_112th_lo;
    end

    // 225. 113th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_113th_hi <= 0;
        else                    reg_64bit_113th_hi <= i_reg_64bit_113th_hi;
    end

    // 226. 113th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_113th_lo <= 0;
        else                    reg_64bit_113th_lo <= i_reg_64bit_113th_lo;
    end

    // 227. 114th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_114th_hi <= 0;
        else                    reg_64bit_114th_hi <= i_reg_64bit_114th_hi;
    end

    // 228. 114th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_114th_lo <= 0;
        else                    reg_64bit_114th_lo <= i_reg_64bit_114th_lo;
    end

    // 229. 115th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_115th_hi <= 0;
        else                    reg_64bit_115th_hi <= i_reg_64bit_115th_hi;
    end

    // 230. 115th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_115th_lo <= 0;
        else                    reg_64bit_115th_lo <= i_reg_64bit_115th_lo;
    end

    // 231. 116th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_116th_hi <= 0;
        else                    reg_64bit_116th_hi <= i_reg_64bit_116th_hi;
    end

    // 232. 116th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_116th_lo <= 0;
        else                    reg_64bit_116th_lo <= i_reg_64bit_116th_lo;
    end

    // 233. 117th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_117th_hi <= 0;
        else                    reg_64bit_117th_hi <= i_reg_64bit_117th_hi;
    end

    // 234. 117th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_117th_lo <= 0;
        else                    reg_64bit_117th_lo <= i_reg_64bit_117th_lo;
    end

    // 235. 118th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_118th_hi <= 0;
        else                    reg_64bit_118th_hi <= i_reg_64bit_118th_hi;
    end

    // 236. 118th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_118th_lo <= 0;
        else                    reg_64bit_118th_lo <= i_reg_64bit_118th_lo;
    end

    // 237. 119th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_119th_hi <= 0;
        else                    reg_64bit_119th_hi <= i_reg_64bit_119th_hi;
    end

    // 238. 119th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_119th_lo <= 0;
        else                    reg_64bit_119th_lo <= i_reg_64bit_119th_lo;
    end

    // 239. 120th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_120th_hi <= 0;
        else                    reg_64bit_120th_hi <= i_reg_64bit_120th_hi;
    end

    // 240. 120th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_120th_lo <= 0;
        else                    reg_64bit_120th_lo <= i_reg_64bit_120th_lo;
    end

    // 241. 121th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_121th_hi <= 0;
        else                    reg_64bit_121th_hi <= i_reg_64bit_121th_hi;
    end

    // 242. 121th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_121th_lo <= 0;
        else                    reg_64bit_121th_lo <= i_reg_64bit_121th_lo;
    end

    // 243. 122th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_122th_hi <= 0;
        else                    reg_64bit_122th_hi <= i_reg_64bit_122th_hi;
    end

    // 244. 122th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_122th_lo <= 0;
        else                    reg_64bit_122th_lo <= i_reg_64bit_122th_lo;
    end

    // 245. 123th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_123th_hi <= 0;
        else                    reg_64bit_123th_hi <= i_reg_64bit_123th_hi;
    end

    // 246. 123th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_123th_lo <= 0;
        else                    reg_64bit_123th_lo <= i_reg_64bit_123th_lo;
    end

    // 247. 124th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_124th_hi <= 0;
        else                    reg_64bit_124th_hi <= i_reg_64bit_124th_hi;
    end

    // 248. 124th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_124th_lo <= 0;
        else                    reg_64bit_124th_lo <= i_reg_64bit_124th_lo;
    end

    // 249. 125th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_125th_hi <= 0;
        else                    reg_64bit_125th_hi <= i_reg_64bit_125th_hi;
    end

    // 250. 125th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_125th_lo <= 0;
        else                    reg_64bit_125th_lo <= i_reg_64bit_125th_lo;
    end

    // 251. 126th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_126th_hi <= 0;
        else                    reg_64bit_126th_hi <= i_reg_64bit_126th_hi;
    end

    // 252. 126th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_126th_lo <= 0;
        else                    reg_64bit_126th_lo <= i_reg_64bit_126th_lo;
    end

    // 253. 127th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_127th_hi <= 0;
        else                    reg_64bit_127th_hi <= i_reg_64bit_127th_hi;
    end

    // 254. 127th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_127th_lo <= 0;
        else                    reg_64bit_127th_lo <= i_reg_64bit_127th_lo;
    end

    // 255. 128th 64-bit Register's Upper Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_128th_hi <= 0;
        else                    reg_64bit_128th_hi <= i_reg_64bit_128th_hi;
    end

    // 256. 128th 64-bit Register's Lower Part
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN)      reg_64bit_128th_lo <= 0;
        else                    reg_64bit_128th_lo <= i_reg_64bit_128th_lo;
    end


// ============================================================================ //
//                                                                              //
//                                  Core Logic                                  //
//                                                                              //
// ============================================================================ //

// ==================================================================== //
//  [1] Comb. Logic for Upper Flag                                      //
// ==================================================================== //
    always @(*) begin
        if(S_AXI_ARVALID & ~S_AXI_ARREADY) begin
            case(S_AXI_ARADDR[OPT_MEM_ADDR_BITS+2:2])
                // # User Guide : Comment the Registers which are Write or Un-Used Registers
                8'h00   :   upper_flag = 1;
                8'h02   :   upper_flag = 1;
                8'h04   :   upper_flag = 1;
                8'h06   :   upper_flag = 1;
                8'h08   :   upper_flag = 1;
                8'h0A   :   upper_flag = 1;
                8'h0C   :   upper_flag = 1;
                8'h0E   :   upper_flag = 1;
                8'h10   :   upper_flag = 1;
                8'h12   :   upper_flag = 1;
                8'h14   :   upper_flag = 1;
                8'h16   :   upper_flag = 1;             
                8'h18   :   upper_flag = 1;
                8'h1A   :   upper_flag = 1;
                8'h1C   :   upper_flag = 1;
                8'h1E   :   upper_flag = 1;
                8'h20   :   upper_flag = 1;
                8'h22   :   upper_flag = 1;
                8'h24   :   upper_flag = 1;
                8'h26   :   upper_flag = 1;
                8'h28   :   upper_flag = 1;
                8'h2A   :   upper_flag = 1;
                8'h2C   :   upper_flag = 1;
                8'h2E   :   upper_flag = 1;
                8'h30   :   upper_flag = 1;
                8'h32   :   upper_flag = 1;
                8'h34   :   upper_flag = 1;
                8'h36   :   upper_flag = 1;
                8'h38   :   upper_flag = 1;
                8'h3A   :   upper_flag = 1;
                8'h3C   :   upper_flag = 1;
                8'h3E   :   upper_flag = 1;
                8'h40   :   upper_flag = 1;
                8'h42   :   upper_flag = 1;
                8'h44   :   upper_flag = 1;
                8'h46   :   upper_flag = 1;
                8'h48   :   upper_flag = 1;
                8'h4A   :   upper_flag = 1;
                8'h4C   :   upper_flag = 1;
                8'h4E   :   upper_flag = 1;
                8'h50   :   upper_flag = 1;
                8'h52   :   upper_flag = 1;
                8'h54   :   upper_flag = 1;
                8'h56   :   upper_flag = 1;
                8'h58   :   upper_flag = 1;
                8'h5A   :   upper_flag = 1;
                8'h5C   :   upper_flag = 1;
                8'h5E   :   upper_flag = 1;
                8'h60   :   upper_flag = 1;
                8'h62   :   upper_flag = 1;
                8'h64   :   upper_flag = 1;
                8'h66   :   upper_flag = 1;
                8'h68   :   upper_flag = 1;
                8'h6A   :   upper_flag = 1;
                8'h6C   :   upper_flag = 1;
                8'h6E   :   upper_flag = 1;
                8'h70   :   upper_flag = 1;
                8'h72   :   upper_flag = 1;
                8'h74   :   upper_flag = 1;
                8'h76   :   upper_flag = 1;
                8'h78   :   upper_flag = 1;
                8'h7A   :   upper_flag = 1;
                8'h7C   :   upper_flag = 1;
                8'h7E   :   upper_flag = 1;
                8'h80   :   upper_flag = 1;
                8'h82   :   upper_flag = 1;
                8'h84   :   upper_flag = 1;
                8'h86   :   upper_flag = 1;
                8'h88   :   upper_flag = 1;
                8'h8A   :   upper_flag = 1;
                8'h8C   :   upper_flag = 1;
                8'h8E   :   upper_flag = 1;
                8'h90   :   upper_flag = 1;
                8'h92   :   upper_flag = 1;
                8'h94   :   upper_flag = 1;
                8'h96   :   upper_flag = 1;
                8'h98   :   upper_flag = 1;
                8'h9A   :   upper_flag = 1;
                8'h9C   :   upper_flag = 1;
                8'h9E   :   upper_flag = 1;
                8'hA0   :   upper_flag = 1;
                8'hA2   :   upper_flag = 1;
                8'hA4   :   upper_flag = 1;
                8'hA6   :   upper_flag = 1;
                8'hA8   :   upper_flag = 1;
                8'hAA   :   upper_flag = 1;
                8'hAC   :   upper_flag = 1;
                8'hAE   :   upper_flag = 1;
                8'hB0   :   upper_flag = 1;
                8'hB2   :   upper_flag = 1;
                8'hB4   :   upper_flag = 1;
                8'hB6   :   upper_flag = 1;
                8'hB8   :   upper_flag = 1;
                8'hBA   :   upper_flag = 1;
                8'hBC   :   upper_flag = 1;
                8'hBE   :   upper_flag = 1;
                8'hC0   :   upper_flag = 1;
                8'hC2   :   upper_flag = 1;
                8'hC4   :   upper_flag = 1;
                8'hC6   :   upper_flag = 1;
                8'hC8   :   upper_flag = 1;
                8'hCA   :   upper_flag = 1;
                8'hCC   :   upper_flag = 1;
                8'hCE   :   upper_flag = 1;
                8'hD0   :   upper_flag = 1;
                8'hD2   :   upper_flag = 1;
                8'hD4   :   upper_flag = 1;
                8'hD6   :   upper_flag = 1;
                8'hD8   :   upper_flag = 1;
                8'hDA   :   upper_flag = 1;
                8'hDC   :   upper_flag = 1;
                8'hDE   :   upper_flag = 1;
                8'hE0   :   upper_flag = 1;
                8'hE2   :   upper_flag = 1;
                8'hE4   :   upper_flag = 1;
                8'hE6   :   upper_flag = 1;
                8'hE8   :   upper_flag = 1;
                8'hEA   :   upper_flag = 1;
                8'hEC   :   upper_flag = 1;
                8'hEE   :   upper_flag = 1;
                8'hF0   :   upper_flag = 1;
                8'hF2   :   upper_flag = 1;
                8'hF4   :   upper_flag = 1;
                8'hF6   :   upper_flag = 1;
                8'hF8   :   upper_flag = 1;
                8'hFA   :   upper_flag = 1;
                8'hFC   :   upper_flag = 1;
                8'hFE   :   upper_flag = 1;
                default :   upper_flag = 0;
            endcase
        end
        else begin
            upper_flag = 0;
        end
    end

// ==================================================================== //
//  [2] Seq. Logic for Register Data Capture                            //
// ==================================================================== //
    always @(posedge S_AXI_ACLK) begin
        if(!S_AXI_ARESETN) begin
            captured_data <= 0;
        end
        else if(upper_flag) begin
            case(S_AXI_ARADDR[OPT_MEM_ADDR_BITS+2:2])
                // # User Guide : Comment the Registers which are Write or Un-Used Registers
                8'h00   :   captured_data <= {reg_64bit_1th_hi, reg_64bit_1th_lo};
                8'h02   :   captured_data <= {reg_64bit_2th_hi, reg_64bit_2th_lo};
                8'h04   :   captured_data <= {reg_64bit_3th_hi, reg_64bit_3th_lo};
                8'h06   :   captured_data <= {reg_64bit_4th_hi, reg_64bit_4th_lo};
                8'h08   :   captured_data <= {reg_64bit_5th_hi, reg_64bit_5th_lo};
                8'h0A   :   captured_data <= {reg_64bit_6th_hi, reg_64bit_6th_lo};
                8'h0C   :   captured_data <= {reg_64bit_7th_hi, reg_64bit_7th_lo};
                8'h0E   :   captured_data <= {reg_64bit_8th_hi, reg_64bit_8th_lo};
                8'h10   :   captured_data <= {reg_64bit_9th_hi, reg_64bit_9th_lo};
                8'h12   :   captured_data <= {reg_64bit_10th_hi, reg_64bit_10th_lo};
                8'h14   :   captured_data <= {reg_64bit_11th_hi, reg_64bit_11th_lo};
                8'h16   :   captured_data <= {reg_64bit_12th_hi, reg_64bit_12th_lo};
                8'h18   :   captured_data <= {reg_64bit_13th_hi, reg_64bit_13th_lo};
                8'h1A   :   captured_data <= {reg_64bit_14th_hi, reg_64bit_14th_lo};
                8'h1C   :   captured_data <= {reg_64bit_15th_hi, reg_64bit_15th_lo};
                8'h1E   :   captured_data <= {reg_64bit_16th_hi, reg_64bit_16th_lo};
                8'h20   :   captured_data <= {reg_64bit_17th_hi, reg_64bit_17th_lo};
                8'h22   :   captured_data <= {reg_64bit_18th_hi, reg_64bit_18th_lo};
                8'h24   :   captured_data <= {reg_64bit_19th_hi, reg_64bit_19th_lo};
                8'h26   :   captured_data <= {reg_64bit_20th_hi, reg_64bit_20th_lo};
                8'h28   :   captured_data <= {reg_64bit_21th_hi, reg_64bit_21th_lo};
                8'h2A   :   captured_data <= {reg_64bit_22th_hi, reg_64bit_22th_lo};
                8'h2C   :   captured_data <= {reg_64bit_23th_hi, reg_64bit_23th_lo};
                8'h2E   :   captured_data <= {reg_64bit_24th_hi, reg_64bit_24th_lo};
                8'h30   :   captured_data <= {reg_64bit_25th_hi, reg_64bit_25th_lo};
                8'h32   :   captured_data <= {reg_64bit_26th_hi, reg_64bit_26th_lo};
                8'h34   :   captured_data <= {reg_64bit_27th_hi, reg_64bit_27th_lo};
                8'h36   :   captured_data <= {reg_64bit_28th_hi, reg_64bit_28th_lo};
                8'h38   :   captured_data <= {reg_64bit_29th_hi, reg_64bit_29th_lo};
                8'h3A   :   captured_data <= {reg_64bit_30th_hi, reg_64bit_30th_lo};
                8'h3C   :   captured_data <= {reg_64bit_31th_hi, reg_64bit_31th_lo};
                8'h3E   :   captured_data <= {reg_64bit_32th_hi, reg_64bit_32th_lo};
                8'h40   :   captured_data <= {reg_64bit_33th_hi, reg_64bit_33th_lo};
                8'h42   :   captured_data <= {reg_64bit_34th_hi, reg_64bit_34th_lo};
                8'h44   :   captured_data <= {reg_64bit_35th_hi, reg_64bit_35th_lo};
                8'h46   :   captured_data <= {reg_64bit_36th_hi, reg_64bit_36th_lo};
                8'h48   :   captured_data <= {reg_64bit_37th_hi, reg_64bit_37th_lo};
                8'h4A   :   captured_data <= {reg_64bit_38th_hi, reg_64bit_38th_lo};
                8'h4C   :   captured_data <= {reg_64bit_39th_hi, reg_64bit_39th_lo};
                8'h4E   :   captured_data <= {reg_64bit_40th_hi, reg_64bit_40th_lo};
                8'h50   :   captured_data <= {reg_64bit_41th_hi, reg_64bit_41th_lo};
                8'h52   :   captured_data <= {reg_64bit_42th_hi, reg_64bit_42th_lo};
                8'h54   :   captured_data <= {reg_64bit_43th_hi, reg_64bit_43th_lo};
                8'h56   :   captured_data <= {reg_64bit_44th_hi, reg_64bit_44th_lo};
                8'h58   :   captured_data <= {reg_64bit_45th_hi, reg_64bit_45th_lo};
                8'h5A   :   captured_data <= {reg_64bit_46th_hi, reg_64bit_46th_lo};
                8'h5C   :   captured_data <= {reg_64bit_47th_hi, reg_64bit_47th_lo};
                8'h5E   :   captured_data <= {reg_64bit_48th_hi, reg_64bit_48th_lo};
                8'h60   :   captured_data <= {reg_64bit_49th_hi, reg_64bit_49th_lo};
                8'h62   :   captured_data <= {reg_64bit_50th_hi, reg_64bit_50th_lo};
                8'h64   :   captured_data <= {reg_64bit_51th_hi, reg_64bit_51th_lo};
                8'h66   :   captured_data <= {reg_64bit_52th_hi, reg_64bit_52th_lo};
                8'h68   :   captured_data <= {reg_64bit_53th_hi, reg_64bit_53th_lo};
                8'h6A   :   captured_data <= {reg_64bit_54th_hi, reg_64bit_54th_lo};
                8'h6C   :   captured_data <= {reg_64bit_55th_hi, reg_64bit_55th_lo};
                8'h6E   :   captured_data <= {reg_64bit_56th_hi, reg_64bit_56th_lo};
                8'h70   :   captured_data <= {reg_64bit_57th_hi, reg_64bit_57th_lo};
                8'h72   :   captured_data <= {reg_64bit_58th_hi, reg_64bit_58th_lo};
                8'h74   :   captured_data <= {reg_64bit_59th_hi, reg_64bit_59th_lo};
                8'h76   :   captured_data <= {reg_64bit_60th_hi, reg_64bit_60th_lo};
                8'h78   :   captured_data <= {reg_64bit_61th_hi, reg_64bit_61th_lo};
                8'h7A   :   captured_data <= {reg_64bit_62th_hi, reg_64bit_62th_lo};
                8'h7C   :   captured_data <= {reg_64bit_63th_hi, reg_64bit_63th_lo};
                8'h7E   :   captured_data <= {reg_64bit_64th_hi, reg_64bit_64th_lo};
                8'h80   :   captured_data <= {reg_64bit_65th_hi, reg_64bit_65th_lo};
                8'h82   :   captured_data <= {reg_64bit_66th_hi, reg_64bit_66th_lo};
                8'h84   :   captured_data <= {reg_64bit_67th_hi, reg_64bit_67th_lo};
                8'h86   :   captured_data <= {reg_64bit_68th_hi, reg_64bit_68th_lo};
                8'h88   :   captured_data <= {reg_64bit_69th_hi, reg_64bit_69th_lo};
                8'h8A   :   captured_data <= {reg_64bit_70th_hi, reg_64bit_70th_lo};
                8'h8C   :   captured_data <= {reg_64bit_71th_hi, reg_64bit_71th_lo};
                8'h8E   :   captured_data <= {reg_64bit_72th_hi, reg_64bit_72th_lo};
                8'h90   :   captured_data <= {reg_64bit_73th_hi, reg_64bit_73th_lo};
                8'h92   :   captured_data <= {reg_64bit_74th_hi, reg_64bit_74th_lo};
                8'h94   :   captured_data <= {reg_64bit_75th_hi, reg_64bit_75th_lo};
                8'h96   :   captured_data <= {reg_64bit_76th_hi, reg_64bit_76th_lo};
                8'h98   :   captured_data <= {reg_64bit_77th_hi, reg_64bit_77th_lo};
                8'h9A   :   captured_data <= {reg_64bit_78th_hi, reg_64bit_78th_lo};
                8'h9C   :   captured_data <= {reg_64bit_79th_hi, reg_64bit_79th_lo};
                8'h9E   :   captured_data <= {reg_64bit_80th_hi, reg_64bit_80th_lo};
                8'hA0   :   captured_data <= {reg_64bit_81th_hi, reg_64bit_81th_lo};
                8'hA2   :   captured_data <= {reg_64bit_82th_hi, reg_64bit_82th_lo};
                8'hA4   :   captured_data <= {reg_64bit_83th_hi, reg_64bit_83th_lo};
                8'hA6   :   captured_data <= {reg_64bit_84th_hi, reg_64bit_84th_lo};
                8'hA8   :   captured_data <= {reg_64bit_85th_hi, reg_64bit_85th_lo};
                8'hAA   :   captured_data <= {reg_64bit_86th_hi, reg_64bit_86th_lo};
                8'hAC   :   captured_data <= {reg_64bit_87th_hi, reg_64bit_87th_lo};
                8'hAE   :   captured_data <= {reg_64bit_88th_hi, reg_64bit_88th_lo};
                8'hB0   :   captured_data <= {reg_64bit_89th_hi, reg_64bit_89th_lo};
                8'hB2   :   captured_data <= {reg_64bit_90th_hi, reg_64bit_90th_lo};
                8'hB4   :   captured_data <= {reg_64bit_91th_hi, reg_64bit_91th_lo};
                8'hB6   :   captured_data <= {reg_64bit_92th_hi, reg_64bit_92th_lo};
                8'hB8   :   captured_data <= {reg_64bit_93th_hi, reg_64bit_93th_lo};
                8'hBA   :   captured_data <= {reg_64bit_94th_hi, reg_64bit_94th_lo};
                8'hBC   :   captured_data <= {reg_64bit_95th_hi, reg_64bit_95th_lo};
                8'hBE   :   captured_data <= {reg_64bit_96th_hi, reg_64bit_96th_lo};
                8'hC0   :   captured_data <= {reg_64bit_97th_hi, reg_64bit_97th_lo};
                8'hC2   :   captured_data <= {reg_64bit_98th_hi, reg_64bit_98th_lo};
                8'hC4   :   captured_data <= {reg_64bit_99th_hi, reg_64bit_99th_lo};
                8'hC6   :   captured_data <= {reg_64bit_100th_hi, reg_64bit_100th_lo};
                8'hC8   :   captured_data <= {reg_64bit_101th_hi, reg_64bit_101th_lo};
                8'hCA   :   captured_data <= {reg_64bit_102th_hi, reg_64bit_102th_lo};
                8'hCC   :   captured_data <= {reg_64bit_103th_hi, reg_64bit_103th_lo};
                8'hCE   :   captured_data <= {reg_64bit_104th_hi, reg_64bit_104th_lo};
                8'hD0   :   captured_data <= {reg_64bit_105th_hi, reg_64bit_105th_lo};
                8'hD2   :   captured_data <= {reg_64bit_106th_hi, reg_64bit_106th_lo};
                8'hD4   :   captured_data <= {reg_64bit_107th_hi, reg_64bit_107th_lo};
                8'hD6   :   captured_data <= {reg_64bit_108th_hi, reg_64bit_108th_lo};
                8'hD8   :   captured_data <= {reg_64bit_109th_hi, reg_64bit_109th_lo};
                8'hDA   :   captured_data <= {reg_64bit_110th_hi, reg_64bit_110th_lo};
                8'hDC   :   captured_data <= {reg_64bit_111th_hi, reg_64bit_111th_lo};
                8'hDE   :   captured_data <= {reg_64bit_112th_hi, reg_64bit_112th_lo};
                8'hE0   :   captured_data <= {reg_64bit_113th_hi, reg_64bit_113th_lo};
                8'hE2   :   captured_data <= {reg_64bit_114th_hi, reg_64bit_114th_lo};
                8'hE4   :   captured_data <= {reg_64bit_115th_hi, reg_64bit_115th_lo};
                8'hE6   :   captured_data <= {reg_64bit_116th_hi, reg_64bit_116th_lo};
                8'hE8   :   captured_data <= {reg_64bit_117th_hi, reg_64bit_117th_lo};
                8'hEA   :   captured_data <= {reg_64bit_118th_hi, reg_64bit_118th_lo};
                8'hEC   :   captured_data <= {reg_64bit_119th_hi, reg_64bit_119th_lo};
                8'hEE   :   captured_data <= {reg_64bit_120th_hi, reg_64bit_120th_lo};
                8'hF0   :   captured_data <= {reg_64bit_121th_hi, reg_64bit_121th_lo};
                8'hF2   :   captured_data <= {reg_64bit_122th_hi, reg_64bit_122th_lo};
                8'hF4   :   captured_data <= {reg_64bit_123th_hi, reg_64bit_123th_lo};
                8'hF6   :   captured_data <= {reg_64bit_124th_hi, reg_64bit_124th_lo};
                8'hF8   :   captured_data <= {reg_64bit_125th_hi, reg_64bit_125th_lo};
                8'hFA   :   captured_data <= {reg_64bit_126th_hi, reg_64bit_126th_lo};
                8'hFC   :   captured_data <= {reg_64bit_127th_hi, reg_64bit_127th_lo};
                8'hFE   :   captured_data <= {reg_64bit_128th_hi, reg_64bit_128th_lo};
                default :   captured_data <= 0;
            endcase
        end
    end

// ==================================================================== //
//  [3] Comb. Logic for Data Source of Slave Registers                  //
// ==================================================================== //
    always @(*) begin
        case(axi_araddr[OPT_MEM_ADDR_BITS+2:2])
            // # User Guide : Comment the Registers which are Write or Un-Used Registers
            8'h00   :   slv_reg0 = captured_data[63:32];
            8'h01   :   slv_reg1 = captured_data[31:0];
            8'h02   :   slv_reg2 = captured_data[63:32];
            8'h03   :   slv_reg3 = captured_data[31:0];
            8'h04   :   slv_reg4 = captured_data[63:32];
            8'h05   :   slv_reg5 = captured_data[31:0];
            8'h06   :   slv_reg6 = captured_data[63:32];
            8'h07   :   slv_reg7 = captured_data[31:0];
            8'h08   :   slv_reg8 = captured_data[63:32];
            8'h09   :   slv_reg9 = captured_data[31:0];
            8'h0A   :   slv_reg10 = captured_data[63:32];
            8'h0B   :   slv_reg11 = captured_data[31:0];
            8'h0C   :   slv_reg12 = captured_data[63:32];
            8'h0D   :   slv_reg13 = captured_data[31:0];
            8'h0E   :   slv_reg14 = captured_data[63:32];
            8'h0F   :   slv_reg15 = captured_data[31:0];
            8'h10   :   slv_reg16 = captured_data[63:32];
            8'h11   :   slv_reg17 = captured_data[31:0];
            8'h12   :   slv_reg18 = captured_data[63:32];
            8'h13   :   slv_reg19 = captured_data[31:0];
            8'h14   :   slv_reg20 = captured_data[63:32];
            8'h15   :   slv_reg21 = captured_data[31:0];
            8'h16   :   slv_reg22 = captured_data[63:32];
            8'h17   :   slv_reg23 = captured_data[31:0];
            8'h18   :   slv_reg24 = captured_data[63:32];
            8'h19   :   slv_reg25 = captured_data[31:0];
            8'h1A   :   slv_reg26 = captured_data[63:32];
            8'h1B   :   slv_reg27 = captured_data[31:0];
            8'h1C   :   slv_reg28 = captured_data[63:32];
            8'h1D   :   slv_reg29 = captured_data[31:0];
            8'h1E   :   slv_reg30 = captured_data[63:32];
            8'h1F   :   slv_reg31 = captured_data[31:0];
            8'h20   :   slv_reg32 = captured_data[63:32];
            8'h21   :   slv_reg33 = captured_data[31:0];
            8'h22   :   slv_reg34 = captured_data[63:32];
            8'h23   :   slv_reg35 = captured_data[31:0];
            8'h24   :   slv_reg36 = captured_data[63:32];
            8'h25   :   slv_reg37 = captured_data[31:0];
            8'h26   :   slv_reg38 = captured_data[63:32];
            8'h27   :   slv_reg39 = captured_data[31:0];
            8'h28   :   slv_reg40 = captured_data[63:32];
            8'h29   :   slv_reg41 = captured_data[31:0];
            8'h2A   :   slv_reg42 = captured_data[63:32];
            8'h2B   :   slv_reg43 = captured_data[31:0];
            8'h2C   :   slv_reg44 = captured_data[63:32];
            8'h2D   :   slv_reg45 = captured_data[31:0];
            8'h2E   :   slv_reg46 = captured_data[63:32];
            8'h2F   :   slv_reg47 = captured_data[31:0];
            8'h30   :   slv_reg48 = captured_data[63:32];
            8'h31   :   slv_reg49 = captured_data[31:0];
            8'h32   :   slv_reg50 = captured_data[63:32];
            8'h33   :   slv_reg51 = captured_data[31:0];
            8'h34   :   slv_reg52 = captured_data[63:32];
            8'h35   :   slv_reg53 = captured_data[31:0];
            8'h36   :   slv_reg54 = captured_data[63:32];
            8'h37   :   slv_reg55 = captured_data[31:0];
            8'h38   :   slv_reg56 = captured_data[63:32];
            8'h39   :   slv_reg57 = captured_data[31:0];
            8'h3A   :   slv_reg58 = captured_data[63:32];
            8'h3B   :   slv_reg59 = captured_data[31:0];
            8'h3C   :   slv_reg60 = captured_data[63:32];
            8'h3D   :   slv_reg61 = captured_data[31:0];
            8'h3E   :   slv_reg62 = captured_data[63:32];
            8'h3F   :   slv_reg63 = captured_data[31:0];
            8'h40   :   slv_reg64 = captured_data[63:32];
            8'h41   :   slv_reg65 = captured_data[31:0];
            8'h42   :   slv_reg66 = captured_data[63:32];
            8'h43   :   slv_reg67 = captured_data[31:0];
            8'h44   :   slv_reg68 = captured_data[63:32];
            8'h45   :   slv_reg69 = captured_data[31:0];
            8'h46   :   slv_reg70 = captured_data[63:32];
            8'h47   :   slv_reg71 = captured_data[31:0];
            8'h48   :   slv_reg72 = captured_data[63:32];
            8'h49   :   slv_reg73 = captured_data[31:0];
            8'h4A   :   slv_reg74 = captured_data[63:32];
            8'h4B   :   slv_reg75 = captured_data[31:0];
            8'h4C   :   slv_reg76 = captured_data[63:32];
            8'h4D   :   slv_reg77 = captured_data[31:0];
            8'h4E   :   slv_reg78 = captured_data[63:32];
            8'h4F   :   slv_reg79 = captured_data[31:0];
            8'h50   :   slv_reg80 = captured_data[63:32];
            8'h51   :   slv_reg81 = captured_data[31:0];
            8'h52   :   slv_reg82 = captured_data[63:32];
            8'h53   :   slv_reg83 = captured_data[31:0];
            8'h54   :   slv_reg84 = captured_data[63:32];
            8'h55   :   slv_reg85 = captured_data[31:0];
            8'h56   :   slv_reg86 = captured_data[63:32];
            8'h57   :   slv_reg87 = captured_data[31:0];
            8'h58   :   slv_reg88 = captured_data[63:32];
            8'h59   :   slv_reg89 = captured_data[31:0];
            8'h5A   :   slv_reg90 = captured_data[63:32];
            8'h5B   :   slv_reg91 = captured_data[31:0];
            8'h5C   :   slv_reg92 = captured_data[63:32];
            8'h5D   :   slv_reg93 = captured_data[31:0];
            8'h5E   :   slv_reg94 = captured_data[63:32];
            8'h5F   :   slv_reg95 = captured_data[31:0];
            8'h60   :   slv_reg96 = captured_data[63:32];
            8'h61   :   slv_reg97 = captured_data[31:0];
            8'h62   :   slv_reg98 = captured_data[63:32];
            8'h63   :   slv_reg99 = captured_data[31:0];
            8'h64   :   slv_reg100 = captured_data[63:32];
            8'h65   :   slv_reg101 = captured_data[31:0];
            8'h66   :   slv_reg102 = captured_data[63:32];
            8'h67   :   slv_reg103 = captured_data[31:0];
            8'h68   :   slv_reg104 = captured_data[63:32];
            8'h69   :   slv_reg105 = captured_data[31:0];
            8'h6A   :   slv_reg106 = captured_data[63:32];
            8'h6B   :   slv_reg107 = captured_data[31:0];
            8'h6C   :   slv_reg108 = captured_data[63:32];
            8'h6D   :   slv_reg109 = captured_data[31:0];
            8'h6E   :   slv_reg110 = captured_data[63:32];
            8'h6F   :   slv_reg111 = captured_data[31:0];
            8'h70   :   slv_reg112 = captured_data[63:32];
            8'h71   :   slv_reg113 = captured_data[31:0];
            8'h72   :   slv_reg114 = captured_data[63:32];
            8'h73   :   slv_reg115 = captured_data[31:0];
            8'h74   :   slv_reg116 = captured_data[63:32];
            8'h75   :   slv_reg117 = captured_data[31:0];
            8'h76   :   slv_reg118 = captured_data[63:32];
            8'h77   :   slv_reg119 = captured_data[31:0];
            8'h78   :   slv_reg120 = captured_data[63:32];
            8'h79   :   slv_reg121 = captured_data[31:0];
            8'h7A   :   slv_reg122 = captured_data[63:32];
            8'h7B   :   slv_reg123 = captured_data[31:0];
            8'h7C   :   slv_reg124 = captured_data[63:32];
            8'h7D   :   slv_reg125 = captured_data[31:0];
            8'h7E   :   slv_reg126 = captured_data[63:32];
            8'h7F   :   slv_reg127 = captured_data[31:0];
            8'h80   :   slv_reg128 = captured_data[63:32];
            8'h81   :   slv_reg129 = captured_data[31:0];
            8'h82   :   slv_reg130 = captured_data[63:32];
            8'h83   :   slv_reg131 = captured_data[31:0];
            8'h84   :   slv_reg132 = captured_data[63:32];
            8'h85   :   slv_reg133 = captured_data[31:0];
            8'h86   :   slv_reg134 = captured_data[63:32];
            8'h87   :   slv_reg135 = captured_data[31:0];
            8'h88   :   slv_reg136 = captured_data[63:32];
            8'h89   :   slv_reg137 = captured_data[31:0];
            8'h8A   :   slv_reg138 = captured_data[63:32];
            8'h8B   :   slv_reg139 = captured_data[31:0];
            8'h8C   :   slv_reg140 = captured_data[63:32];
            8'h8D   :   slv_reg141 = captured_data[31:0];
            8'h8E   :   slv_reg142 = captured_data[63:32];
            8'h8F   :   slv_reg143 = captured_data[31:0];
            8'h90   :   slv_reg144 = captured_data[63:32];
            8'h91   :   slv_reg145 = captured_data[31:0];
            8'h92   :   slv_reg146 = captured_data[63:32];
            8'h93   :   slv_reg147 = captured_data[31:0];
            8'h94   :   slv_reg148 = captured_data[63:32];
            8'h95   :   slv_reg149 = captured_data[31:0];
            8'h96   :   slv_reg150 = captured_data[63:32];
            8'h97   :   slv_reg151 = captured_data[31:0];
            8'h98   :   slv_reg152 = captured_data[63:32];
            8'h99   :   slv_reg153 = captured_data[31:0];
            8'h9A   :   slv_reg154 = captured_data[63:32];
            8'h9B   :   slv_reg155 = captured_data[31:0];
            8'h9C   :   slv_reg156 = captured_data[63:32];
            8'h9D   :   slv_reg157 = captured_data[31:0];
            8'h9E   :   slv_reg158 = captured_data[63:32];
            8'h9F   :   slv_reg159 = captured_data[31:0];
            8'hA0   :   slv_reg160 = captured_data[63:32];
            8'hA1   :   slv_reg161 = captured_data[31:0];
            8'hA2   :   slv_reg162 = captured_data[63:32];
            8'hA3   :   slv_reg163 = captured_data[31:0];
            8'hA4   :   slv_reg164 = captured_data[63:32];
            8'hA5   :   slv_reg165 = captured_data[31:0];
            8'hA6   :   slv_reg166 = captured_data[63:32];
            8'hA7   :   slv_reg167 = captured_data[31:0];
            8'hA8   :   slv_reg168 = captured_data[63:32];
            8'hA9   :   slv_reg169 = captured_data[31:0];
            8'hAA   :   slv_reg170 = captured_data[63:32];
            8'hAB   :   slv_reg171 = captured_data[31:0];
            8'hAC   :   slv_reg172 = captured_data[63:32];
            8'hAD   :   slv_reg173 = captured_data[31:0];
            8'hAE   :   slv_reg174 = captured_data[63:32];
            8'hAF   :   slv_reg175 = captured_data[31:0];
            8'hB0   :   slv_reg176 = captured_data[63:32];
            8'hB1   :   slv_reg177 = captured_data[31:0];
            8'hB2   :   slv_reg178 = captured_data[63:32];
            8'hB3   :   slv_reg179 = captured_data[31:0];
            8'hB4   :   slv_reg180 = captured_data[63:32];
            8'hB5   :   slv_reg181 = captured_data[31:0];
            8'hB6   :   slv_reg182 = captured_data[63:32];
            8'hB7   :   slv_reg183 = captured_data[31:0];
            8'hB8   :   slv_reg184 = captured_data[63:32];
            8'hB9   :   slv_reg185 = captured_data[31:0];
            8'hBA   :   slv_reg186 = captured_data[63:32];
            8'hBB   :   slv_reg187 = captured_data[31:0];
            8'hBC   :   slv_reg188 = captured_data[63:32];
            8'hBD   :   slv_reg189 = captured_data[31:0];
            8'hBE   :   slv_reg190 = captured_data[63:32];
            8'hBF   :   slv_reg191 = captured_data[31:0];
            8'hC0   :   slv_reg192 = captured_data[63:32];
            8'hC1   :   slv_reg193 = captured_data[31:0];
            8'hC2   :   slv_reg194 = captured_data[63:32];
            8'hC3   :   slv_reg195 = captured_data[31:0];
            8'hC4   :   slv_reg196 = captured_data[63:32];
            8'hC5   :   slv_reg197 = captured_data[31:0];
            8'hC6   :   slv_reg198 = captured_data[63:32];
            8'hC7   :   slv_reg199 = captured_data[31:0];
            8'hC8   :   slv_reg200 = captured_data[63:32];
            8'hC9   :   slv_reg201 = captured_data[31:0];
            8'hCA   :   slv_reg202 = captured_data[63:32];
            8'hCB   :   slv_reg203 = captured_data[31:0];
            8'hCC   :   slv_reg204 = captured_data[63:32];
            8'hCD   :   slv_reg205 = captured_data[31:0];
            8'hCE   :   slv_reg206 = captured_data[63:32];
            8'hCF   :   slv_reg207 = captured_data[31:0];
            8'hD0   :   slv_reg208 = captured_data[63:32];
            8'hD1   :   slv_reg209 = captured_data[31:0];
            8'hD2   :   slv_reg210 = captured_data[63:32];
            8'hD3   :   slv_reg211 = captured_data[31:0];
            8'hD4   :   slv_reg212 = captured_data[63:32];
            8'hD5   :   slv_reg213 = captured_data[31:0];
            8'hD6   :   slv_reg214 = captured_data[63:32];
            8'hD7   :   slv_reg215 = captured_data[31:0];
            8'hD8   :   slv_reg216 = captured_data[63:32];
            8'hD9   :   slv_reg217 = captured_data[31:0];
            8'hDA   :   slv_reg218 = captured_data[63:32];
            8'hDB   :   slv_reg219 = captured_data[31:0];
            8'hDC   :   slv_reg220 = captured_data[63:32];
            8'hDD   :   slv_reg221 = captured_data[31:0];
            8'hDE   :   slv_reg222 = captured_data[63:32];
            8'hDF   :   slv_reg223 = captured_data[31:0];
            8'hE0   :   slv_reg224 = captured_data[63:32];
            8'hE1   :   slv_reg225 = captured_data[31:0];
            8'hE2   :   slv_reg226 = captured_data[63:32];
            8'hE3   :   slv_reg227 = captured_data[31:0];
            8'hE4   :   slv_reg228 = captured_data[63:32];
            8'hE5   :   slv_reg229 = captured_data[31:0];
            8'hE6   :   slv_reg230 = captured_data[63:32];
            8'hE7   :   slv_reg231 = captured_data[31:0];
            8'hE8   :   slv_reg232 = captured_data[63:32];
            8'hE9   :   slv_reg233 = captured_data[31:0];
            8'hEA   :   slv_reg234 = captured_data[63:32];
            8'hEB   :   slv_reg235 = captured_data[31:0];
            8'hEC   :   slv_reg236 = captured_data[63:32];
            8'hED   :   slv_reg237 = captured_data[31:0];
            8'hEE   :   slv_reg238 = captured_data[63:32];
            8'hEF   :   slv_reg239 = captured_data[31:0];
            8'hF0   :   slv_reg240 = captured_data[63:32];
            8'hF1   :   slv_reg241 = captured_data[31:0];
            8'hF2   :   slv_reg242 = captured_data[63:32];
            8'hF3   :   slv_reg243 = captured_data[31:0];
            8'hF4   :   slv_reg244 = captured_data[63:32];
            8'hF5   :   slv_reg245 = captured_data[31:0];
            8'hF6   :   slv_reg246 = captured_data[63:32];
            8'hF7   :   slv_reg247 = captured_data[31:0];
            8'hF8   :   slv_reg248 = captured_data[63:32];
            8'hF9   :   slv_reg249 = captured_data[31:0];
            8'hFA   :   slv_reg250 = captured_data[63:32];
            8'hFB   :   slv_reg251 = captured_data[31:0];
            8'hFC   :   slv_reg252 = captured_data[63:32];
            8'hFD   :   slv_reg253 = captured_data[31:0];
            8'hFE   :   slv_reg254 = captured_data[63:32];
            8'hFF   :   slv_reg255 = captured_data[31:0];
            default : begin
                        // # User Guide : Comment the Registers which are Write or Un-Used Registers
                        slv_reg0 = 0;
                        slv_reg1 = 0;
                        slv_reg2 = 0;
                        slv_reg3 = 0;
                        slv_reg4 = 0;
                        slv_reg5 = 0;
                        slv_reg6 = 0;
                        slv_reg7 = 0;
                        slv_reg8 = 0;
                        slv_reg9 = 0;
                        slv_reg10 = 0;
                        slv_reg11 = 0;
                        slv_reg12 = 0;
                        slv_reg13 = 0;
                        slv_reg14 = 0;
                        slv_reg15 = 0;
                        slv_reg16 = 0;
                        slv_reg17 = 0;
                        slv_reg18 = 0;
                        slv_reg19 = 0;
                        slv_reg20 = 0;
                        slv_reg21 = 0;
                        slv_reg22 = 0;
                        slv_reg23 = 0;
                        slv_reg24 = 0;
                        slv_reg25 = 0;
                        slv_reg26 = 0;
                        slv_reg27 = 0;
                        slv_reg28 = 0;
                        slv_reg29 = 0;
                        slv_reg30 = 0;
                        slv_reg31 = 0;
                        slv_reg32 = 0;
                        slv_reg33 = 0;
                        slv_reg34 = 0;
                        slv_reg35 = 0;
                        slv_reg36 = 0;
                        slv_reg37 = 0;
                        slv_reg38 = 0;
                        slv_reg39 = 0;
                        slv_reg40 = 0;
                        slv_reg41 = 0;
                        slv_reg42 = 0;
                        slv_reg43 = 0;
                        slv_reg44 = 0;
                        slv_reg45 = 0;
                        slv_reg46 = 0;
                        slv_reg47 = 0;
                        slv_reg48 = 0;
                        slv_reg49 = 0;
                        slv_reg50 = 0;
                        slv_reg51 = 0;
                        slv_reg52 = 0;
                        slv_reg53 = 0;
                        slv_reg54 = 0;
                        slv_reg55 = 0;
                        slv_reg56 = 0;
                        slv_reg57 = 0;
                        slv_reg58 = 0;
                        slv_reg59 = 0;
                        slv_reg60 = 0;
                        slv_reg61 = 0;
                        slv_reg62 = 0;
                        slv_reg63 = 0;
                        slv_reg64 = 0;
                        slv_reg65 = 0;
                        slv_reg66 = 0;
                        slv_reg67 = 0;
                        slv_reg68 = 0;
                        slv_reg69 = 0;
                        slv_reg70 = 0;
                        slv_reg71 = 0;
                        slv_reg72 = 0;
                        slv_reg73 = 0;
                        slv_reg74 = 0;
                        slv_reg75 = 0;
                        slv_reg76 = 0;
                        slv_reg77 = 0;
                        slv_reg78 = 0;
                        slv_reg79 = 0;
                        slv_reg80 = 0;
                        slv_reg81 = 0;
                        slv_reg82 = 0;
                        slv_reg83 = 0;
                        slv_reg84 = 0;
                        slv_reg85 = 0;
                        slv_reg86 = 0;
                        slv_reg87 = 0;
                        slv_reg88 = 0;
                        slv_reg89 = 0;
                        slv_reg90 = 0;
                        slv_reg91 = 0;
                        slv_reg92 = 0;
                        slv_reg93 = 0;
                        slv_reg94 = 0;
                        slv_reg95 = 0;
                        slv_reg96 = 0;
                        slv_reg97 = 0;
                        slv_reg98 = 0;
                        slv_reg99 = 0;
                        slv_reg100 = 0;
                        slv_reg101 = 0;
                        slv_reg102 = 0;
                        slv_reg103 = 0;
                        slv_reg104 = 0;
                        slv_reg105 = 0;
                        slv_reg106 = 0;
                        slv_reg107 = 0;
                        slv_reg108 = 0;
                        slv_reg109 = 0;
                        slv_reg110 = 0;
                        slv_reg111 = 0;
                        slv_reg112 = 0;
                        slv_reg113 = 0;
                        slv_reg114 = 0;
                        slv_reg115 = 0;
                        slv_reg116 = 0;
                        slv_reg117 = 0;
                        slv_reg118 = 0;
                        slv_reg119 = 0;
                        slv_reg120 = 0;
                        slv_reg121 = 0;
                        slv_reg122 = 0;
                        slv_reg123 = 0;
                        slv_reg124 = 0;
                        slv_reg125 = 0;
                        slv_reg126 = 0;
                        slv_reg127 = 0;
                        slv_reg128 = 0;
                        slv_reg129 = 0;
                        slv_reg130 = 0;
                        slv_reg131 = 0;
                        slv_reg132 = 0;
                        slv_reg133 = 0;
                        slv_reg134 = 0;
                        slv_reg135 = 0;
                        slv_reg136 = 0;
                        slv_reg137 = 0;
                        slv_reg138 = 0;
                        slv_reg139 = 0;
                        slv_reg140 = 0;
                        slv_reg141 = 0;
                        slv_reg142 = 0;
                        slv_reg143 = 0;
                        slv_reg144 = 0;
                        slv_reg145 = 0;
                        slv_reg146 = 0;
                        slv_reg147 = 0;
                        slv_reg148 = 0;
                        slv_reg149 = 0;
                        slv_reg150 = 0;
                        slv_reg151 = 0;
                        slv_reg152 = 0;
                        slv_reg153 = 0;
                        slv_reg154 = 0;
                        slv_reg155 = 0;
                        slv_reg156 = 0;
                        slv_reg157 = 0;
                        slv_reg158 = 0;
                        slv_reg159 = 0;
                        slv_reg160 = 0;
                        slv_reg161 = 0;
                        slv_reg162 = 0;
                        slv_reg163 = 0;
                        slv_reg164 = 0;
                        slv_reg165 = 0;
                        slv_reg166 = 0;
                        slv_reg167 = 0;
                        slv_reg168 = 0;
                        slv_reg169 = 0;
                        slv_reg170 = 0;
                        slv_reg171 = 0;
                        slv_reg172 = 0;
                        slv_reg173 = 0;
                        slv_reg174 = 0;
                        slv_reg175 = 0;
                        slv_reg176 = 0;
                        slv_reg177 = 0;
                        slv_reg178 = 0;
                        slv_reg179 = 0;
                        slv_reg180 = 0;
                        slv_reg181 = 0;
                        slv_reg182 = 0;
                        slv_reg183 = 0;
                        slv_reg184 = 0;
                        slv_reg185 = 0;
                        slv_reg186 = 0;
                        slv_reg187 = 0;
                        slv_reg188 = 0;
                        slv_reg189 = 0;
                        slv_reg190 = 0;
                        slv_reg191 = 0;
                        slv_reg192 = 0;
                        slv_reg193 = 0;
                        slv_reg194 = 0;
                        slv_reg195 = 0;
                        slv_reg196 = 0;
                        slv_reg197 = 0;
                        slv_reg198 = 0;
                        slv_reg199 = 0;
                        slv_reg200 = 0;
                        slv_reg201 = 0;
                        slv_reg202 = 0;
                        slv_reg203 = 0;
                        slv_reg204 = 0;
                        slv_reg205 = 0;
                        slv_reg206 = 0;
                        slv_reg207 = 0;
                        slv_reg208 = 0;
                        slv_reg209 = 0;
                        slv_reg210 = 0;
                        slv_reg211 = 0;
                        slv_reg212 = 0;
                        slv_reg213 = 0;
                        slv_reg214 = 0;
                        slv_reg215 = 0;
                        slv_reg216 = 0;
                        slv_reg217 = 0;
                        slv_reg218 = 0;
                        slv_reg219 = 0;
                        slv_reg220 = 0;
                        slv_reg221 = 0;
                        slv_reg222 = 0;
                        slv_reg223 = 0;
                        slv_reg224 = 0;
                        slv_reg225 = 0;
                        slv_reg226 = 0;
                        slv_reg227 = 0;
                        slv_reg228 = 0;
                        slv_reg229 = 0;
                        slv_reg230 = 0;
                        slv_reg231 = 0;
                        slv_reg232 = 0;
                        slv_reg233 = 0;
                        slv_reg234 = 0;
                        slv_reg235 = 0;
                        slv_reg236 = 0;
                        slv_reg237 = 0;
                        slv_reg238 = 0;
                        slv_reg239 = 0;
                        slv_reg240 = 0;
                        slv_reg241 = 0;
                        slv_reg242 = 0;
                        slv_reg243 = 0;
                        slv_reg244 = 0;
                        slv_reg245 = 0;
                        slv_reg246 = 0;
                        slv_reg247 = 0;
                        slv_reg248 = 0;
                        slv_reg249 = 0;
                        slv_reg250 = 0;
                        slv_reg251 = 0;
                        slv_reg252 = 0;
                        slv_reg253 = 0;
                        slv_reg254 = 0;
                        slv_reg255 = 0;
                    end
        endcase
    end


// ============================================================================ //
//                                                                              //
//                              Output Assignments                              //
//                                                                              //
// ============================================================================ //
    // # User Guide : Un-Comment the Pins which are Connected to Write Registers
    // assign  o_reg_64bit_1th_hi = slv_reg0;
    // assign  o_reg_64bit_1th_lo = slv_reg1;
    // assign  o_reg_64bit_2th_hi = slv_reg2;
    // assign  o_reg_64bit_2th_lo = slv_reg3;
    // assign  o_reg_64bit_3th_hi = slv_reg4;
    // assign  o_reg_64bit_3th_lo = slv_reg5;
    // assign  o_reg_64bit_4th_hi = slv_reg6;
    // assign  o_reg_64bit_4th_lo = slv_reg7;
    // assign  o_reg_64bit_5th_hi = slv_reg8;
    // assign  o_reg_64bit_5th_lo = slv_reg9;
    // assign  o_reg_64bit_6th_hi = slv_reg10;
    // assign  o_reg_64bit_6th_lo = slv_reg11;
    // assign  o_reg_64bit_7th_hi = slv_reg12;
    // assign  o_reg_64bit_7th_lo = slv_reg13;
    // assign  o_reg_64bit_8th_hi = slv_reg14;
    // assign  o_reg_64bit_8th_lo = slv_reg15;
    // assign  o_reg_64bit_9th_hi = slv_reg16;
    // assign  o_reg_64bit_9th_lo = slv_reg17;
    // assign  o_reg_64bit_10th_hi = slv_reg18;
    // assign  o_reg_64bit_10th_lo = slv_reg19;
    // assign  o_reg_64bit_11th_hi = slv_reg20;
    // assign  o_reg_64bit_11th_lo = slv_reg21;
    // assign  o_reg_64bit_12th_hi = slv_reg22;
    // assign  o_reg_64bit_12th_lo = slv_reg23;
    // assign  o_reg_64bit_13th_hi = slv_reg24;
    // assign  o_reg_64bit_13th_lo = slv_reg25;
    // assign  o_reg_64bit_14th_hi = slv_reg26;
    // assign  o_reg_64bit_14th_lo = slv_reg27;
    // assign  o_reg_64bit_15th_hi = slv_reg28;
    // assign  o_reg_64bit_15th_lo = slv_reg29;
    // assign  o_reg_64bit_16th_hi = slv_reg30;
    // assign  o_reg_64bit_16th_lo = slv_reg31;
    // assign  o_reg_64bit_17th_hi = slv_reg32;
    // assign  o_reg_64bit_17th_lo = slv_reg33;
    // assign  o_reg_64bit_18th_hi = slv_reg34;
    // assign  o_reg_64bit_18th_lo = slv_reg35;
    // assign  o_reg_64bit_19th_hi = slv_reg36;
    // assign  o_reg_64bit_19th_lo = slv_reg37;
    // assign  o_reg_64bit_20th_hi = slv_reg38;
    // assign  o_reg_64bit_20th_lo = slv_reg39;
    // assign  o_reg_64bit_21th_hi = slv_reg40;
    // assign  o_reg_64bit_21th_lo = slv_reg41;
    // assign  o_reg_64bit_22th_hi = slv_reg42;
    // assign  o_reg_64bit_22th_lo = slv_reg43;
    // assign  o_reg_64bit_23th_hi = slv_reg44;
    // assign  o_reg_64bit_23th_lo = slv_reg45;
    // assign  o_reg_64bit_24th_hi = slv_reg46;
    // assign  o_reg_64bit_24th_lo = slv_reg47;
    // assign  o_reg_64bit_25th_hi = slv_reg48;
    // assign  o_reg_64bit_25th_lo = slv_reg49;
    // assign  o_reg_64bit_26th_hi = slv_reg50;
    // assign  o_reg_64bit_26th_lo = slv_reg51;
    // assign  o_reg_64bit_27th_hi = slv_reg52;
    // assign  o_reg_64bit_27th_lo = slv_reg53;
    // assign  o_reg_64bit_28th_hi = slv_reg54;
    // assign  o_reg_64bit_28th_lo = slv_reg55;
    // assign  o_reg_64bit_29th_hi = slv_reg56;
    // assign  o_reg_64bit_29th_lo = slv_reg57;
    // assign  o_reg_64bit_30th_hi = slv_reg58;
    // assign  o_reg_64bit_30th_lo = slv_reg59;
    // assign  o_reg_64bit_31th_hi = slv_reg60;
    // assign  o_reg_64bit_31th_lo = slv_reg61;
    // assign  o_reg_64bit_32th_hi = slv_reg62;
    // assign  o_reg_64bit_32th_lo = slv_reg63;
    // assign  o_reg_64bit_33th_hi = slv_reg64;
    // assign  o_reg_64bit_33th_lo = slv_reg65;
    // assign  o_reg_64bit_34th_hi = slv_reg66;
    // assign  o_reg_64bit_34th_lo = slv_reg67;
    // assign  o_reg_64bit_35th_hi = slv_reg68;
    // assign  o_reg_64bit_35th_lo = slv_reg69;
    // assign  o_reg_64bit_36th_hi = slv_reg70;
    // assign  o_reg_64bit_36th_lo = slv_reg71;
    // assign  o_reg_64bit_37th_hi = slv_reg72;
    // assign  o_reg_64bit_37th_lo = slv_reg73;
    // assign  o_reg_64bit_38th_hi = slv_reg74;
    // assign  o_reg_64bit_38th_lo = slv_reg75;
    // assign  o_reg_64bit_39th_hi = slv_reg76;
    // assign  o_reg_64bit_39th_lo = slv_reg77;
    // assign  o_reg_64bit_40th_hi = slv_reg78;
    // assign  o_reg_64bit_40th_lo = slv_reg79;
    // assign  o_reg_64bit_41th_hi = slv_reg80;
    // assign  o_reg_64bit_41th_lo = slv_reg81;
    // assign  o_reg_64bit_42th_hi = slv_reg82;
    // assign  o_reg_64bit_42th_lo = slv_reg83;
    // assign  o_reg_64bit_43th_hi = slv_reg84;
    // assign  o_reg_64bit_43th_lo = slv_reg85;
    // assign  o_reg_64bit_44th_hi = slv_reg86;
    // assign  o_reg_64bit_44th_lo = slv_reg87;
    // assign  o_reg_64bit_45th_hi = slv_reg88;
    // assign  o_reg_64bit_45th_lo = slv_reg89;
    // assign  o_reg_64bit_46th_hi = slv_reg90;
    // assign  o_reg_64bit_46th_lo = slv_reg91;
    // assign  o_reg_64bit_47th_hi = slv_reg92;
    // assign  o_reg_64bit_47th_lo = slv_reg93;
    // assign  o_reg_64bit_48th_hi = slv_reg94;
    // assign  o_reg_64bit_48th_lo = slv_reg95;
    // assign  o_reg_64bit_49th_hi = slv_reg96;
    // assign  o_reg_64bit_49th_lo = slv_reg97;
    // assign  o_reg_64bit_50th_hi = slv_reg98;
    // assign  o_reg_64bit_50th_lo = slv_reg99;
    // assign  o_reg_64bit_51th_hi = slv_reg100;
    // assign  o_reg_64bit_51th_lo = slv_reg101;
    // assign  o_reg_64bit_52th_hi = slv_reg102;
    // assign  o_reg_64bit_52th_lo = slv_reg103;
    // assign  o_reg_64bit_53th_hi = slv_reg104;
    // assign  o_reg_64bit_53th_lo = slv_reg105;
    // assign  o_reg_64bit_54th_hi = slv_reg106;
    // assign  o_reg_64bit_54th_lo = slv_reg107;
    // assign  o_reg_64bit_55th_hi = slv_reg108;
    // assign  o_reg_64bit_55th_lo = slv_reg109;
    // assign  o_reg_64bit_56th_hi = slv_reg110;
    // assign  o_reg_64bit_56th_lo = slv_reg111;
    // assign  o_reg_64bit_57th_hi = slv_reg112;
    // assign  o_reg_64bit_57th_lo = slv_reg113;
    // assign  o_reg_64bit_58th_hi = slv_reg114;
    // assign  o_reg_64bit_58th_lo = slv_reg115;
    // assign  o_reg_64bit_59th_hi = slv_reg116;
    // assign  o_reg_64bit_59th_lo = slv_reg117;
    // assign  o_reg_64bit_60th_hi = slv_reg118;
    // assign  o_reg_64bit_60th_lo = slv_reg119;
    // assign  o_reg_64bit_61th_hi = slv_reg120;
    // assign  o_reg_64bit_61th_lo = slv_reg121;
    // assign  o_reg_64bit_62th_hi = slv_reg122;
    // assign  o_reg_64bit_62th_lo = slv_reg123;
    // assign  o_reg_64bit_63th_hi = slv_reg124;
    // assign  o_reg_64bit_63th_lo = slv_reg125;
    // assign  o_reg_64bit_64th_hi = slv_reg126;
    // assign  o_reg_64bit_64th_lo = slv_reg127;
    // assign  o_reg_64bit_65th_hi = slv_reg128;
    // assign  o_reg_64bit_65th_lo = slv_reg129;
    // assign  o_reg_64bit_66th_hi = slv_reg130;
    // assign  o_reg_64bit_66th_lo = slv_reg131;
    // assign  o_reg_64bit_67th_hi = slv_reg132;
    // assign  o_reg_64bit_67th_lo = slv_reg133;
    // assign  o_reg_64bit_68th_hi = slv_reg134;
    // assign  o_reg_64bit_68th_lo = slv_reg135;
    // assign  o_reg_64bit_69th_hi = slv_reg136;
    // assign  o_reg_64bit_69th_lo = slv_reg137;
    // assign  o_reg_64bit_70th_hi = slv_reg138;
    // assign  o_reg_64bit_70th_lo = slv_reg139;
    // assign  o_reg_64bit_71th_hi = slv_reg140;
    // assign  o_reg_64bit_71th_lo = slv_reg141;
    // assign  o_reg_64bit_72th_hi = slv_reg142;
    // assign  o_reg_64bit_72th_lo = slv_reg143;
    // assign  o_reg_64bit_73th_hi = slv_reg144;
    // assign  o_reg_64bit_73th_lo = slv_reg145;
    // assign  o_reg_64bit_74th_hi = slv_reg146;
    // assign  o_reg_64bit_74th_lo = slv_reg147;
    // assign  o_reg_64bit_75th_hi = slv_reg148;
    // assign  o_reg_64bit_75th_lo = slv_reg149;
    // assign  o_reg_64bit_76th_hi = slv_reg150;
    // assign  o_reg_64bit_76th_lo = slv_reg151;
    // assign  o_reg_64bit_77th_hi = slv_reg152;
    // assign  o_reg_64bit_77th_lo = slv_reg153;
    // assign  o_reg_64bit_78th_hi = slv_reg154;
    // assign  o_reg_64bit_78th_lo = slv_reg155;
    // assign  o_reg_64bit_79th_hi = slv_reg156;
    // assign  o_reg_64bit_79th_lo = slv_reg157;
    // assign  o_reg_64bit_80th_hi = slv_reg158;
    // assign  o_reg_64bit_80th_lo = slv_reg159;
    // assign  o_reg_64bit_81th_hi = slv_reg160;
    // assign  o_reg_64bit_81th_lo = slv_reg161;
    // assign  o_reg_64bit_82th_hi = slv_reg162;
    // assign  o_reg_64bit_82th_lo = slv_reg163;
    // assign  o_reg_64bit_83th_hi = slv_reg164;
    // assign  o_reg_64bit_83th_lo = slv_reg165;
    // assign  o_reg_64bit_84th_hi = slv_reg166;
    // assign  o_reg_64bit_84th_lo = slv_reg167;
    // assign  o_reg_64bit_85th_hi = slv_reg168;
    // assign  o_reg_64bit_85th_lo = slv_reg169;
    // assign  o_reg_64bit_86th_hi = slv_reg170;
    // assign  o_reg_64bit_86th_lo = slv_reg171;
    // assign  o_reg_64bit_87th_hi = slv_reg172;
    // assign  o_reg_64bit_87th_lo = slv_reg173;
    // assign  o_reg_64bit_88th_hi = slv_reg174;
    // assign  o_reg_64bit_88th_lo = slv_reg175;
    // assign  o_reg_64bit_89th_hi = slv_reg176;
    // assign  o_reg_64bit_89th_lo = slv_reg177;
    // assign  o_reg_64bit_90th_hi = slv_reg178;
    // assign  o_reg_64bit_90th_lo = slv_reg179;
    // assign  o_reg_64bit_91th_hi = slv_reg180;
    // assign  o_reg_64bit_91th_lo = slv_reg181;
    // assign  o_reg_64bit_92th_hi = slv_reg182;
    // assign  o_reg_64bit_92th_lo = slv_reg183;
    // assign  o_reg_64bit_93th_hi = slv_reg184;
    // assign  o_reg_64bit_93th_lo = slv_reg185;
    // assign  o_reg_64bit_94th_hi = slv_reg186;
    // assign  o_reg_64bit_94th_lo = slv_reg187;
    // assign  o_reg_64bit_95th_hi = slv_reg188;
    // assign  o_reg_64bit_95th_lo = slv_reg189;
    // assign  o_reg_64bit_96th_hi = slv_reg190;
    // assign  o_reg_64bit_96th_lo = slv_reg191;
    // assign  o_reg_64bit_97th_hi = slv_reg192;
    // assign  o_reg_64bit_97th_lo = slv_reg193;
    // assign  o_reg_64bit_98th_hi = slv_reg194;
    // assign  o_reg_64bit_98th_lo = slv_reg195;
    // assign  o_reg_64bit_99th_hi = slv_reg196;
    // assign  o_reg_64bit_99th_lo = slv_reg197;
    // assign  o_reg_64bit_100th_hi = slv_reg198;
    // assign  o_reg_64bit_100th_lo = slv_reg199;
    // assign  o_reg_64bit_101th_hi = slv_reg200;
    // assign  o_reg_64bit_101th_lo = slv_reg201;
    // assign  o_reg_64bit_102th_hi = slv_reg202;
    // assign  o_reg_64bit_102th_lo = slv_reg203;
    // assign  o_reg_64bit_103th_hi = slv_reg204;
    // assign  o_reg_64bit_103th_lo = slv_reg205;
    // assign  o_reg_64bit_104th_hi = slv_reg206;
    // assign  o_reg_64bit_104th_lo = slv_reg207;
    // assign  o_reg_64bit_105th_hi = slv_reg208;
    // assign  o_reg_64bit_105th_lo = slv_reg209;
    // assign  o_reg_64bit_106th_hi = slv_reg210;
    // assign  o_reg_64bit_106th_lo = slv_reg211;
    // assign  o_reg_64bit_107th_hi = slv_reg212;
    // assign  o_reg_64bit_107th_lo = slv_reg213;
    // assign  o_reg_64bit_108th_hi = slv_reg214;
    // assign  o_reg_64bit_108th_lo = slv_reg215;
    // assign  o_reg_64bit_109th_hi = slv_reg216;
    // assign  o_reg_64bit_109th_lo = slv_reg217;
    // assign  o_reg_64bit_110th_hi = slv_reg218;
    // assign  o_reg_64bit_110th_lo = slv_reg219;
    // assign  o_reg_64bit_111th_hi = slv_reg220;
    // assign  o_reg_64bit_111th_lo = slv_reg221;
    // assign  o_reg_64bit_112th_hi = slv_reg222;
    // assign  o_reg_64bit_112th_lo = slv_reg223;
    // assign  o_reg_64bit_113th_hi = slv_reg224;
    // assign  o_reg_64bit_113th_lo = slv_reg225;
    // assign  o_reg_64bit_114th_hi = slv_reg226;
    // assign  o_reg_64bit_114th_lo = slv_reg227;
    // assign  o_reg_64bit_115th_hi = slv_reg228;
    // assign  o_reg_64bit_115th_lo = slv_reg229;
    // assign  o_reg_64bit_116th_hi = slv_reg230;
    // assign  o_reg_64bit_116th_lo = slv_reg231;
    // assign  o_reg_64bit_117th_hi = slv_reg232;
    // assign  o_reg_64bit_117th_lo = slv_reg233;
    // assign  o_reg_64bit_118th_hi = slv_reg234;
    // assign  o_reg_64bit_118th_lo = slv_reg235;
    // assign  o_reg_64bit_119th_hi = slv_reg236;
    // assign  o_reg_64bit_119th_lo = slv_reg237;
    // assign  o_reg_64bit_120th_hi = slv_reg238;
    // assign  o_reg_64bit_120th_lo = slv_reg239;
    // assign  o_reg_64bit_121th_hi = slv_reg240;
    // assign  o_reg_64bit_121th_lo = slv_reg241;
    // assign  o_reg_64bit_122th_hi = slv_reg242;
    // assign  o_reg_64bit_122th_lo = slv_reg243;
    // assign  o_reg_64bit_123th_hi = slv_reg244;
    // assign  o_reg_64bit_123th_lo = slv_reg245;
    // assign  o_reg_64bit_124th_hi = slv_reg246;
    // assign  o_reg_64bit_124th_lo = slv_reg247;
    // assign  o_reg_64bit_125th_hi = slv_reg248;
    // assign  o_reg_64bit_125th_lo = slv_reg249;
    // assign  o_reg_64bit_126th_hi = slv_reg250;
    // assign  o_reg_64bit_126th_lo = slv_reg251;
    // assign  o_reg_64bit_127th_hi = slv_reg252;
    // assign  o_reg_64bit_127th_lo = slv_reg253;
    // assign  o_reg_64bit_128th_hi = slv_reg254;
    // assign  o_reg_64bit_128th_lo = slv_reg255;

endmodule
